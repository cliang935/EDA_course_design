`timescale 1ns/10ps

module wtree_4to2_64x64(
  input    wire        clk  ,
  input    wire        rstn ,
  input    wire [65:0] pp1  ,
  input    wire [65:0] pp2  ,
  input    wire [65:0] pp3  ,
  input    wire [65:0] pp4  ,
  input    wire [65:0] pp5  ,
  input    wire [65:0] pp6  ,
  input    wire [65:0] pp7  ,
  input    wire [65:0] pp8  ,
  input    wire [65:0] pp9  ,
  input    wire [65:0] pp10 ,
  input    wire [65:0] pp11 ,
  input    wire [65:0] pp12 ,
  input    wire [65:0] pp13 ,
  input    wire [65:0] pp14 ,
  input    wire [65:0] pp15 ,
  input    wire [65:0] pp16 ,
  input    wire [65:0] pp17 ,
  input    wire [65:0] pp18 ,
  input    wire [65:0] pp19 ,
  input    wire [65:0] pp20 ,
  input    wire [65:0] pp21 ,
  input    wire [65:0] pp22 ,
  input    wire [65:0] pp23 ,
  input    wire [65:0] pp24 ,
  input    wire [65:0] pp25 ,
  input    wire [65:0] pp26 ,
  input    wire [65:0] pp27 ,
  input    wire [65:0] pp28 ,
  input    wire [65:0] pp29 ,
  input    wire [65:0] pp30 ,
  input    wire [65:0] pp31 ,
  input    wire [65:0] pp32 ,
  input    wire [65:0] pp33 ,
  output   wire [127:0] final_p
);

// ================ first stage ================
wire [65:0] pp1_w;
wire [65:0] pp2_w;
wire [65:0] pp3_w;
wire [65:0] pp4_w;
wire [65:0] pp5_w;
wire [65:0] pp6_w;
wire [65:0] pp7_w;
wire [65:0] pp8_w;
wire [65:0] pp9_w;
wire [65:0] pp10_w;
wire [65:0] pp11_w;
wire [65:0] pp12_w;
wire [65:0] pp13_w;
wire [65:0] pp14_w;
wire [65:0] pp15_w;
wire [65:0] pp16_w;
wire [65:0] pp17_w;
wire [65:0] pp18_w;
wire [65:0] pp19_w;
wire [65:0] pp20_w;
wire [65:0] pp21_w;
wire [65:0] pp22_w;
wire [65:0] pp23_w;
wire [65:0] pp24_w;
wire [65:0] pp25_w;
wire [65:0] pp26_w;
wire [65:0] pp27_w;
wire [65:0] pp28_w;
wire [65:0] pp29_w;
wire [65:0] pp30_w;
wire [65:0] pp31_w;
wire [65:0] pp32_w;
wire [65:0] pp33_w;

// ============== pipeline ===============
reg [65:0] pp1_ff ;
reg [65:0] pp2_ff ;
reg [65:0] pp3_ff ;
reg [65:0] pp4_ff ;
reg [65:0] pp5_ff ;
reg [65:0] pp6_ff ;
reg [65:0] pp7_ff ;
reg [65:0] pp8_ff ;
reg [65:0] pp9_ff ;
reg [65:0] pp10_ff;
reg [65:0] pp11_ff;
reg [65:0] pp12_ff;
reg [65:0] pp13_ff;
reg [65:0] pp14_ff;
reg [65:0] pp15_ff;
reg [65:0] pp16_ff;
reg [65:0] pp17_ff;
reg [65:0] pp18_ff;
reg [65:0] pp19_ff;
reg [65:0] pp20_ff;
reg [65:0] pp21_ff;
reg [65:0] pp22_ff;
reg [65:0] pp23_ff;
reg [65:0] pp24_ff;
reg [65:0] pp25_ff;
reg [65:0] pp26_ff;
reg [65:0] pp27_ff;
reg [65:0] pp28_ff;
reg [65:0] pp29_ff;
reg [65:0] pp30_ff;
reg [65:0] pp31_ff;
reg [65:0] pp32_ff;
reg [65:0] pp33_ff;

always @(posedge clk or negedge rstn)begin
    if (!rstn)begin
        pp1_ff  <= 66'b0;
        pp2_ff  <= 66'b0;
        pp3_ff  <= 66'b0;
        pp4_ff  <= 66'b0;
        pp5_ff  <= 66'b0;
        pp6_ff  <= 66'b0;
        pp7_ff  <= 66'b0;
        pp8_ff  <= 66'b0;
        pp9_ff  <= 66'b0;
        pp10_ff <= 66'b0;
        pp11_ff <= 66'b0;
        pp12_ff <= 66'b0;
        pp13_ff <= 66'b0;
        pp14_ff <= 66'b0;
        pp15_ff <= 66'b0;
        pp16_ff <= 66'b0;
        pp17_ff <= 66'b0;
        pp18_ff <= 66'b0;
        pp19_ff <= 66'b0;
        pp20_ff <= 66'b0;
        pp21_ff <= 66'b0;
        pp22_ff <= 66'b0;
        pp23_ff <= 66'b0;
        pp24_ff <= 66'b0;
        pp25_ff <= 66'b0;
        pp26_ff <= 66'b0;
        pp27_ff <= 66'b0;
        pp28_ff <= 66'b0;
        pp29_ff <= 66'b0;
        pp30_ff <= 66'b0;
        pp31_ff <= 66'b0;
        pp32_ff <= 66'b0;
        pp33_ff <= 66'b0;
    end
    else begin
        pp1_ff  <= pp1  ;
        pp2_ff  <= pp2  ;
        pp3_ff  <= pp3  ;
        pp4_ff  <= pp4  ;
        pp5_ff  <= pp5  ;
        pp6_ff  <= pp6  ;
        pp7_ff  <= pp7  ;
        pp8_ff  <= pp8  ;
        pp9_ff  <= pp9  ;
        pp10_ff <= pp10 ;
        pp11_ff <= pp11 ;
        pp12_ff <= pp12 ;
        pp13_ff <= pp13 ;
        pp14_ff <= pp14 ;
        pp15_ff <= pp15 ;
        pp16_ff <= pp16 ;
        pp17_ff <= pp17 ;
        pp18_ff <= pp18 ;
        pp19_ff <= pp19 ;
        pp20_ff <= pp20 ;
        pp21_ff <= pp21 ;
        pp22_ff <= pp22 ;
        pp23_ff <= pp23 ;
        pp24_ff <= pp24 ;
        pp25_ff <= pp25 ;
        pp26_ff <= pp26 ;
        pp27_ff <= pp27 ;
        pp28_ff <= pp28 ;
        pp29_ff <= pp29 ;
        pp30_ff <= pp30 ;
        pp31_ff <= pp31 ;
        pp32_ff <= pp32 ;
        pp33_ff <= pp33 ;
    end
end

assign pp1_w  = pp1_ff  ;
assign pp2_w  = pp2_ff  ;
assign pp3_w  = pp3_ff  ;
assign pp4_w  = pp4_ff  ;
assign pp5_w  = pp5_ff  ;
assign pp6_w  = pp6_ff  ;
assign pp7_w  = pp7_ff  ;
assign pp8_w  = pp8_ff  ;
assign pp9_w  = pp9_ff  ;
assign pp10_w = pp10_ff ;
assign pp11_w = pp11_ff ;
assign pp12_w = pp12_ff ;
assign pp13_w = pp13_ff ;
assign pp14_w = pp14_ff ;
assign pp15_w = pp15_ff ;
assign pp16_w = pp16_ff ;
assign pp17_w = pp17_ff ;
assign pp18_w = pp18_ff ;
assign pp19_w = pp19_ff ;
assign pp20_w = pp20_ff ;
assign pp21_w = pp21_ff ;
assign pp22_w = pp22_ff ;
assign pp23_w = pp23_ff ;
assign pp24_w = pp24_ff ;
assign pp25_w = pp25_ff ;
assign pp26_w = pp26_ff ;
assign pp27_w = pp27_ff ;
assign pp28_w = pp28_ff ;
assign pp29_w = pp29_ff ;
assign pp30_w = pp30_ff ;
assign pp31_w = pp31_ff ;
assign pp32_w = pp32_ff ;
assign pp33_w = pp33_ff ;

wire [72:0] stg1_s1, stg1_c1, stg1_co1;
wire [72:0] stg1_s2, stg1_c2, stg1_co2;
wire [72:0] stg1_s3, stg1_c3, stg1_co3;
wire [72:0] stg1_s4, stg1_c4, stg1_co4;
wire [72:0] stg1_s5, stg1_c5, stg1_co5;
wire [72:0] stg1_s6, stg1_c6, stg1_co6;
wire [72:0] stg1_s7, stg1_c7, stg1_co7;
wire [71:0] stg1_s8, stg1_c8, stg1_co8;

// =========================== first stage 1st group ============================================================================================================
counter_5to3 u_a11_0 (.i0(pp1_w[0 ]), .i1(1'b0     ), .i2(1'b0     ), .i3(1'b0     ), .ci(1'b0        ), .s(stg1_s1[0 ]), .c(stg1_c1[0 ]), .co(stg1_co1[0 ]));
counter_5to3 u_a11_1 (.i0(pp1_w[1 ]), .i1(1'b0     ), .i2(1'b0     ), .i3(1'b0     ), .ci(stg1_co1[0 ]), .s(stg1_s1[1 ]), .c(stg1_c1[1 ]), .co(stg1_co1[1 ]));
counter_5to3 u_a11_2 (.i0(pp1_w[2 ]), .i1(pp2_w[0 ]), .i2(1'b0     ), .i3(1'b0     ), .ci(stg1_co1[1 ]), .s(stg1_s1[2 ]), .c(stg1_c1[2 ]), .co(stg1_co1[2 ]));
counter_5to3 u_a11_3 (.i0(pp1_w[3 ]), .i1(pp2_w[1 ]), .i2(1'b0     ), .i3(1'b0     ), .ci(stg1_co1[2 ]), .s(stg1_s1[3 ]), .c(stg1_c1[3 ]), .co(stg1_co1[3 ]));
counter_5to3 u_a11_4 (.i0(pp1_w[4 ]), .i1(pp2_w[2 ]), .i2(pp3_w[0 ]), .i3(1'b0     ), .ci(stg1_co1[3 ]), .s(stg1_s1[4 ]), .c(stg1_c1[4 ]), .co(stg1_co1[4 ]));
counter_5to3 u_a11_5 (.i0(pp1_w[5 ]), .i1(pp2_w[3 ]), .i2(pp3_w[1 ]), .i3(1'b0     ), .ci(stg1_co1[4 ]), .s(stg1_s1[5 ]), .c(stg1_c1[5 ]), .co(stg1_co1[5 ]));
counter_5to3 u_a11_6 (.i0(pp1_w[6 ]), .i1(pp2_w[4 ]), .i2(pp3_w[2 ]), .i3(pp4_w[0 ]), .ci(stg1_co1[5 ]), .s(stg1_s1[6 ]), .c(stg1_c1[6 ]), .co(stg1_co1[6 ]));
counter_5to3 u_a11_7 (.i0(pp1_w[7 ]), .i1(pp2_w[5 ]), .i2(pp3_w[3 ]), .i3(pp4_w[1 ]), .ci(stg1_co1[6 ]), .s(stg1_s1[7 ]), .c(stg1_c1[7 ]), .co(stg1_co1[7 ]));
counter_5to3 u_a11_8 (.i0(pp1_w[8 ]), .i1(pp2_w[6 ]), .i2(pp3_w[4 ]), .i3(pp4_w[2 ]), .ci(stg1_co1[7 ]), .s(stg1_s1[8 ]), .c(stg1_c1[8 ]), .co(stg1_co1[8 ]));
counter_5to3 u_a11_9 (.i0(pp1_w[9 ]), .i1(pp2_w[7 ]), .i2(pp3_w[5 ]), .i3(pp4_w[3 ]), .ci(stg1_co1[8 ]), .s(stg1_s1[9 ]), .c(stg1_c1[9 ]), .co(stg1_co1[9 ]));
counter_5to3 u_a11_10(.i0(pp1_w[10]), .i1(pp2_w[8 ]), .i2(pp3_w[6 ]), .i3(pp4_w[4 ]), .ci(stg1_co1[9 ]), .s(stg1_s1[10]), .c(stg1_c1[10]), .co(stg1_co1[10]));
counter_5to3 u_a11_11(.i0(pp1_w[11]), .i1(pp2_w[9 ]), .i2(pp3_w[7 ]), .i3(pp4_w[5 ]), .ci(stg1_co1[10]), .s(stg1_s1[11]), .c(stg1_c1[11]), .co(stg1_co1[11]));
counter_5to3 u_a11_12(.i0(pp1_w[12]), .i1(pp2_w[10]), .i2(pp3_w[8 ]), .i3(pp4_w[6 ]), .ci(stg1_co1[11]), .s(stg1_s1[12]), .c(stg1_c1[12]), .co(stg1_co1[12]));
counter_5to3 u_a11_13(.i0(pp1_w[13]), .i1(pp2_w[11]), .i2(pp3_w[9 ]), .i3(pp4_w[7 ]), .ci(stg1_co1[12]), .s(stg1_s1[13]), .c(stg1_c1[13]), .co(stg1_co1[13]));
counter_5to3 u_a11_14(.i0(pp1_w[14]), .i1(pp2_w[12]), .i2(pp3_w[10]), .i3(pp4_w[8 ]), .ci(stg1_co1[13]), .s(stg1_s1[14]), .c(stg1_c1[14]), .co(stg1_co1[14]));
counter_5to3 u_a11_15(.i0(pp1_w[15]), .i1(pp2_w[13]), .i2(pp3_w[11]), .i3(pp4_w[9 ]), .ci(stg1_co1[14]), .s(stg1_s1[15]), .c(stg1_c1[15]), .co(stg1_co1[15]));
counter_5to3 u_a11_16(.i0(pp1_w[16]), .i1(pp2_w[14]), .i2(pp3_w[12]), .i3(pp4_w[10]), .ci(stg1_co1[15]), .s(stg1_s1[16]), .c(stg1_c1[16]), .co(stg1_co1[16]));
counter_5to3 u_a11_17(.i0(pp1_w[17]), .i1(pp2_w[15]), .i2(pp3_w[13]), .i3(pp4_w[11]), .ci(stg1_co1[16]), .s(stg1_s1[17]), .c(stg1_c1[17]), .co(stg1_co1[17]));
counter_5to3 u_a11_18(.i0(pp1_w[18]), .i1(pp2_w[16]), .i2(pp3_w[14]), .i3(pp4_w[12]), .ci(stg1_co1[17]), .s(stg1_s1[18]), .c(stg1_c1[18]), .co(stg1_co1[18]));
counter_5to3 u_a11_19(.i0(pp1_w[19]), .i1(pp2_w[17]), .i2(pp3_w[15]), .i3(pp4_w[13]), .ci(stg1_co1[18]), .s(stg1_s1[19]), .c(stg1_c1[19]), .co(stg1_co1[19]));
counter_5to3 u_a11_20(.i0(pp1_w[20]), .i1(pp2_w[18]), .i2(pp3_w[16]), .i3(pp4_w[14]), .ci(stg1_co1[19]), .s(stg1_s1[20]), .c(stg1_c1[20]), .co(stg1_co1[20]));
counter_5to3 u_a11_21(.i0(pp1_w[21]), .i1(pp2_w[19]), .i2(pp3_w[17]), .i3(pp4_w[15]), .ci(stg1_co1[20]), .s(stg1_s1[21]), .c(stg1_c1[21]), .co(stg1_co1[21]));
counter_5to3 u_a11_22(.i0(pp1_w[22]), .i1(pp2_w[20]), .i2(pp3_w[18]), .i3(pp4_w[16]), .ci(stg1_co1[21]), .s(stg1_s1[22]), .c(stg1_c1[22]), .co(stg1_co1[22]));
counter_5to3 u_a11_23(.i0(pp1_w[23]), .i1(pp2_w[21]), .i2(pp3_w[19]), .i3(pp4_w[17]), .ci(stg1_co1[22]), .s(stg1_s1[23]), .c(stg1_c1[23]), .co(stg1_co1[23]));
counter_5to3 u_a11_24(.i0(pp1_w[24]), .i1(pp2_w[22]), .i2(pp3_w[20]), .i3(pp4_w[18]), .ci(stg1_co1[23]), .s(stg1_s1[24]), .c(stg1_c1[24]), .co(stg1_co1[24]));
counter_5to3 u_a11_25(.i0(pp1_w[25]), .i1(pp2_w[23]), .i2(pp3_w[21]), .i3(pp4_w[19]), .ci(stg1_co1[24]), .s(stg1_s1[25]), .c(stg1_c1[25]), .co(stg1_co1[25]));
counter_5to3 u_a11_26(.i0(pp1_w[26]), .i1(pp2_w[24]), .i2(pp3_w[22]), .i3(pp4_w[20]), .ci(stg1_co1[25]), .s(stg1_s1[26]), .c(stg1_c1[26]), .co(stg1_co1[26]));
counter_5to3 u_a11_27(.i0(pp1_w[27]), .i1(pp2_w[25]), .i2(pp3_w[23]), .i3(pp4_w[21]), .ci(stg1_co1[26]), .s(stg1_s1[27]), .c(stg1_c1[27]), .co(stg1_co1[27]));
counter_5to3 u_a11_28(.i0(pp1_w[28]), .i1(pp2_w[26]), .i2(pp3_w[24]), .i3(pp4_w[22]), .ci(stg1_co1[27]), .s(stg1_s1[28]), .c(stg1_c1[28]), .co(stg1_co1[28]));
counter_5to3 u_a11_29(.i0(pp1_w[29]), .i1(pp2_w[27]), .i2(pp3_w[25]), .i3(pp4_w[23]), .ci(stg1_co1[28]), .s(stg1_s1[29]), .c(stg1_c1[29]), .co(stg1_co1[29]));
counter_5to3 u_a11_30(.i0(pp1_w[30]), .i1(pp2_w[28]), .i2(pp3_w[26]), .i3(pp4_w[24]), .ci(stg1_co1[29]), .s(stg1_s1[30]), .c(stg1_c1[30]), .co(stg1_co1[30]));
counter_5to3 u_a11_31(.i0(pp1_w[31]), .i1(pp2_w[29]), .i2(pp3_w[27]), .i3(pp4_w[25]), .ci(stg1_co1[30]), .s(stg1_s1[31]), .c(stg1_c1[31]), .co(stg1_co1[31]));
counter_5to3 u_a11_32(.i0(pp1_w[32]), .i1(pp2_w[30]), .i2(pp3_w[28]), .i3(pp4_w[26]), .ci(stg1_co1[31]), .s(stg1_s1[32]), .c(stg1_c1[32]), .co(stg1_co1[32]));
counter_5to3 u_a11_33(.i0(pp1_w[33]), .i1(pp2_w[31]), .i2(pp3_w[29]), .i3(pp4_w[27]), .ci(stg1_co1[32]), .s(stg1_s1[33]), .c(stg1_c1[33]), .co(stg1_co1[33]));
counter_5to3 u_a11_34(.i0(pp1_w[34]), .i1(pp2_w[32]), .i2(pp3_w[30]), .i3(pp4_w[28]), .ci(stg1_co1[33]), .s(stg1_s1[34]), .c(stg1_c1[34]), .co(stg1_co1[34]));
counter_5to3 u_a11_35(.i0(pp1_w[35]), .i1(pp2_w[33]), .i2(pp3_w[31]), .i3(pp4_w[29]), .ci(stg1_co1[34]), .s(stg1_s1[35]), .c(stg1_c1[35]), .co(stg1_co1[35]));
counter_5to3 u_a11_36(.i0(pp1_w[36]), .i1(pp2_w[34]), .i2(pp3_w[32]), .i3(pp4_w[30]), .ci(stg1_co1[35]), .s(stg1_s1[36]), .c(stg1_c1[36]), .co(stg1_co1[36]));
counter_5to3 u_a11_37(.i0(pp1_w[37]), .i1(pp2_w[35]), .i2(pp3_w[33]), .i3(pp4_w[31]), .ci(stg1_co1[36]), .s(stg1_s1[37]), .c(stg1_c1[37]), .co(stg1_co1[37]));
counter_5to3 u_a11_38(.i0(pp1_w[38]), .i1(pp2_w[36]), .i2(pp3_w[34]), .i3(pp4_w[32]), .ci(stg1_co1[37]), .s(stg1_s1[38]), .c(stg1_c1[38]), .co(stg1_co1[38]));
counter_5to3 u_a11_39(.i0(pp1_w[39]), .i1(pp2_w[37]), .i2(pp3_w[35]), .i3(pp4_w[33]), .ci(stg1_co1[38]), .s(stg1_s1[39]), .c(stg1_c1[39]), .co(stg1_co1[39]));
counter_5to3 u_a11_40(.i0(pp1_w[40]), .i1(pp2_w[38]), .i2(pp3_w[36]), .i3(pp4_w[34]), .ci(stg1_co1[39]), .s(stg1_s1[40]), .c(stg1_c1[40]), .co(stg1_co1[40]));
counter_5to3 u_a11_41(.i0(pp1_w[41]), .i1(pp2_w[39]), .i2(pp3_w[37]), .i3(pp4_w[35]), .ci(stg1_co1[40]), .s(stg1_s1[41]), .c(stg1_c1[41]), .co(stg1_co1[41]));
counter_5to3 u_a11_42(.i0(pp1_w[42]), .i1(pp2_w[40]), .i2(pp3_w[38]), .i3(pp4_w[36]), .ci(stg1_co1[41]), .s(stg1_s1[42]), .c(stg1_c1[42]), .co(stg1_co1[42]));
counter_5to3 u_a11_43(.i0(pp1_w[43]), .i1(pp2_w[41]), .i2(pp3_w[39]), .i3(pp4_w[37]), .ci(stg1_co1[42]), .s(stg1_s1[43]), .c(stg1_c1[43]), .co(stg1_co1[43]));
counter_5to3 u_a11_44(.i0(pp1_w[44]), .i1(pp2_w[42]), .i2(pp3_w[40]), .i3(pp4_w[38]), .ci(stg1_co1[43]), .s(stg1_s1[44]), .c(stg1_c1[44]), .co(stg1_co1[44]));
counter_5to3 u_a11_45(.i0(pp1_w[45]), .i1(pp2_w[43]), .i2(pp3_w[41]), .i3(pp4_w[39]), .ci(stg1_co1[44]), .s(stg1_s1[45]), .c(stg1_c1[45]), .co(stg1_co1[45]));
counter_5to3 u_a11_46(.i0(pp1_w[46]), .i1(pp2_w[44]), .i2(pp3_w[42]), .i3(pp4_w[40]), .ci(stg1_co1[45]), .s(stg1_s1[46]), .c(stg1_c1[46]), .co(stg1_co1[46]));
counter_5to3 u_a11_47(.i0(pp1_w[47]), .i1(pp2_w[45]), .i2(pp3_w[43]), .i3(pp4_w[41]), .ci(stg1_co1[46]), .s(stg1_s1[47]), .c(stg1_c1[47]), .co(stg1_co1[47]));
counter_5to3 u_a11_48(.i0(pp1_w[48]), .i1(pp2_w[46]), .i2(pp3_w[44]), .i3(pp4_w[42]), .ci(stg1_co1[47]), .s(stg1_s1[48]), .c(stg1_c1[48]), .co(stg1_co1[48]));
counter_5to3 u_a11_49(.i0(pp1_w[49]), .i1(pp2_w[47]), .i2(pp3_w[45]), .i3(pp4_w[43]), .ci(stg1_co1[48]), .s(stg1_s1[49]), .c(stg1_c1[49]), .co(stg1_co1[49]));
counter_5to3 u_a11_50(.i0(pp1_w[50]), .i1(pp2_w[48]), .i2(pp3_w[46]), .i3(pp4_w[44]), .ci(stg1_co1[49]), .s(stg1_s1[50]), .c(stg1_c1[50]), .co(stg1_co1[50]));
counter_5to3 u_a11_51(.i0(pp1_w[51]), .i1(pp2_w[49]), .i2(pp3_w[47]), .i3(pp4_w[45]), .ci(stg1_co1[50]), .s(stg1_s1[51]), .c(stg1_c1[51]), .co(stg1_co1[51]));
counter_5to3 u_a11_52(.i0(pp1_w[52]), .i1(pp2_w[50]), .i2(pp3_w[48]), .i3(pp4_w[46]), .ci(stg1_co1[51]), .s(stg1_s1[52]), .c(stg1_c1[52]), .co(stg1_co1[52]));
counter_5to3 u_a11_53(.i0(pp1_w[53]), .i1(pp2_w[51]), .i2(pp3_w[49]), .i3(pp4_w[47]), .ci(stg1_co1[52]), .s(stg1_s1[53]), .c(stg1_c1[53]), .co(stg1_co1[53]));
counter_5to3 u_a11_54(.i0(pp1_w[54]), .i1(pp2_w[52]), .i2(pp3_w[50]), .i3(pp4_w[48]), .ci(stg1_co1[53]), .s(stg1_s1[54]), .c(stg1_c1[54]), .co(stg1_co1[54]));
counter_5to3 u_a11_55(.i0(pp1_w[55]), .i1(pp2_w[53]), .i2(pp3_w[51]), .i3(pp4_w[49]), .ci(stg1_co1[54]), .s(stg1_s1[55]), .c(stg1_c1[55]), .co(stg1_co1[55]));
counter_5to3 u_a11_56(.i0(pp1_w[56]), .i1(pp2_w[54]), .i2(pp3_w[52]), .i3(pp4_w[50]), .ci(stg1_co1[55]), .s(stg1_s1[56]), .c(stg1_c1[56]), .co(stg1_co1[56]));
counter_5to3 u_a11_57(.i0(pp1_w[57]), .i1(pp2_w[55]), .i2(pp3_w[53]), .i3(pp4_w[51]), .ci(stg1_co1[56]), .s(stg1_s1[57]), .c(stg1_c1[57]), .co(stg1_co1[57]));
counter_5to3 u_a11_58(.i0(pp1_w[58]), .i1(pp2_w[56]), .i2(pp3_w[54]), .i3(pp4_w[52]), .ci(stg1_co1[57]), .s(stg1_s1[58]), .c(stg1_c1[58]), .co(stg1_co1[58]));
counter_5to3 u_a11_59(.i0(pp1_w[59]), .i1(pp2_w[57]), .i2(pp3_w[55]), .i3(pp4_w[53]), .ci(stg1_co1[58]), .s(stg1_s1[59]), .c(stg1_c1[59]), .co(stg1_co1[59]));
counter_5to3 u_a11_60(.i0(pp1_w[60]), .i1(pp2_w[58]), .i2(pp3_w[56]), .i3(pp4_w[54]), .ci(stg1_co1[59]), .s(stg1_s1[60]), .c(stg1_c1[60]), .co(stg1_co1[60]));
counter_5to3 u_a11_61(.i0(pp1_w[61]), .i1(pp2_w[59]), .i2(pp3_w[57]), .i3(pp4_w[55]), .ci(stg1_co1[60]), .s(stg1_s1[61]), .c(stg1_c1[61]), .co(stg1_co1[61]));
counter_5to3 u_a11_62(.i0(pp1_w[62]), .i1(pp2_w[60]), .i2(pp3_w[58]), .i3(pp4_w[56]), .ci(stg1_co1[61]), .s(stg1_s1[62]), .c(stg1_c1[62]), .co(stg1_co1[62]));
counter_5to3 u_a11_63(.i0(pp1_w[63]), .i1(pp2_w[61]), .i2(pp3_w[59]), .i3(pp4_w[57]), .ci(stg1_co1[62]), .s(stg1_s1[63]), .c(stg1_c1[63]), .co(stg1_co1[63]));
counter_5to3 u_a11_64(.i0(pp1_w[64]), .i1(pp2_w[62]), .i2(pp3_w[60]), .i3(pp4_w[58]), .ci(stg1_co1[63]), .s(stg1_s1[64]), .c(stg1_c1[64]), .co(stg1_co1[64]));
counter_5to3 u_a11_65(.i0(pp1_w[65]), .i1(pp2_w[63]), .i2(pp3_w[61]), .i3(pp4_w[59]), .ci(stg1_co1[64]), .s(stg1_s1[65]), .c(stg1_c1[65]), .co(stg1_co1[65]));
counter_5to3 u_a11_66(.i0(pp1_w[65]), .i1(pp2_w[64]), .i2(pp3_w[62]), .i3(pp4_w[60]), .ci(stg1_co1[65]), .s(stg1_s1[66]), .c(stg1_c1[66]), .co(stg1_co1[66]));
counter_5to3 u_a11_67(.i0(pp1_w[65]), .i1(pp2_w[65]), .i2(pp3_w[63]), .i3(pp4_w[61]), .ci(stg1_co1[66]), .s(stg1_s1[67]), .c(stg1_c1[67]), .co(stg1_co1[67]));
counter_5to3 u_a11_68(.i0(pp1_w[65]), .i1(pp2_w[65]), .i2(pp3_w[64]), .i3(pp4_w[62]), .ci(stg1_co1[67]), .s(stg1_s1[68]), .c(stg1_c1[68]), .co(stg1_co1[68]));
counter_5to3 u_a11_69(.i0(pp1_w[65]), .i1(pp2_w[65]), .i2(pp3_w[65]), .i3(pp4_w[63]), .ci(stg1_co1[68]), .s(stg1_s1[69]), .c(stg1_c1[69]), .co(stg1_co1[69]));
counter_5to3 u_a11_70(.i0(pp1_w[65]), .i1(pp2_w[65]), .i2(pp3_w[65]), .i3(pp4_w[64]), .ci(stg1_co1[69]), .s(stg1_s1[70]), .c(stg1_c1[70]), .co(stg1_co1[70]));
counter_5to3 u_all_71(.i0(pp1_w[65]), .i1(pp2_w[65]), .i2(pp3_w[65]), .i3(pp4_w[65]), .ci(stg1_co1[70]), .s(stg1_s1[71]), .c(stg1_c1[71]), .co(stg1_co1[71]));
counter_5to3 u_all_72(.i0(pp1_w[65]), .i1(pp2_w[65]), .i2(pp3_w[65]), .i3(pp4_w[65]), .ci(stg1_co1[71]), .s(stg1_s1[72]), .c(stg1_c1[72]), .co(stg1_co1[72]));

// =========================== first stage 2nd group ============================================================================================================
counter_5to3 u_a12_0 (.i0(pp5_w[0 ]), .i1(1'b0     ), .i2(1'b0     ), .i3(1'b0     ), .ci(1'b0        ), .s(stg1_s2[0 ]), .c(stg1_c2[0 ]), .co(stg1_co2[0 ]));
counter_5to3 u_a12_1 (.i0(pp5_w[1 ]), .i1(1'b0     ), .i2(1'b0     ), .i3(1'b0     ), .ci(stg1_co2[0 ]), .s(stg1_s2[1 ]), .c(stg1_c2[1 ]), .co(stg1_co2[1 ]));
counter_5to3 u_a12_2 (.i0(pp5_w[2 ]), .i1(pp6_w[0 ]), .i2(1'b0     ), .i3(1'b0     ), .ci(stg1_co2[1 ]), .s(stg1_s2[2 ]), .c(stg1_c2[2 ]), .co(stg1_co2[2 ]));
counter_5to3 u_a12_3 (.i0(pp5_w[3 ]), .i1(pp6_w[1 ]), .i2(1'b0     ), .i3(1'b0     ), .ci(stg1_co2[2 ]), .s(stg1_s2[3 ]), .c(stg1_c2[3 ]), .co(stg1_co2[3 ]));
counter_5to3 u_a12_4 (.i0(pp5_w[4 ]), .i1(pp6_w[2 ]), .i2(pp7_w[0 ]), .i3(1'b0     ), .ci(stg1_co2[3 ]), .s(stg1_s2[4 ]), .c(stg1_c2[4 ]), .co(stg1_co2[4 ]));
counter_5to3 u_a12_5 (.i0(pp5_w[5 ]), .i1(pp6_w[3 ]), .i2(pp7_w[1 ]), .i3(1'b0     ), .ci(stg1_co2[4 ]), .s(stg1_s2[5 ]), .c(stg1_c2[5 ]), .co(stg1_co2[5 ]));
counter_5to3 u_a12_6 (.i0(pp5_w[6 ]), .i1(pp6_w[4 ]), .i2(pp7_w[2 ]), .i3(pp8_w[0 ]), .ci(stg1_co2[5 ]), .s(stg1_s2[6 ]), .c(stg1_c2[6 ]), .co(stg1_co2[6 ]));
counter_5to3 u_a12_7 (.i0(pp5_w[7 ]), .i1(pp6_w[5 ]), .i2(pp7_w[3 ]), .i3(pp8_w[1 ]), .ci(stg1_co2[6 ]), .s(stg1_s2[7 ]), .c(stg1_c2[7 ]), .co(stg1_co2[7 ]));
counter_5to3 u_a12_8 (.i0(pp5_w[8 ]), .i1(pp6_w[6 ]), .i2(pp7_w[4 ]), .i3(pp8_w[2 ]), .ci(stg1_co2[7 ]), .s(stg1_s2[8 ]), .c(stg1_c2[8 ]), .co(stg1_co2[8 ]));
counter_5to3 u_a12_9 (.i0(pp5_w[9 ]), .i1(pp6_w[7 ]), .i2(pp7_w[5 ]), .i3(pp8_w[3 ]), .ci(stg1_co2[8 ]), .s(stg1_s2[9 ]), .c(stg1_c2[9 ]), .co(stg1_co2[9 ]));
counter_5to3 u_a12_10(.i0(pp5_w[10]), .i1(pp6_w[8 ]), .i2(pp7_w[6 ]), .i3(pp8_w[4 ]), .ci(stg1_co2[9 ]), .s(stg1_s2[10]), .c(stg1_c2[10]), .co(stg1_co2[10]));
counter_5to3 u_a12_11(.i0(pp5_w[11]), .i1(pp6_w[9 ]), .i2(pp7_w[7 ]), .i3(pp8_w[5 ]), .ci(stg1_co2[10]), .s(stg1_s2[11]), .c(stg1_c2[11]), .co(stg1_co2[11]));
counter_5to3 u_a12_12(.i0(pp5_w[12]), .i1(pp6_w[10]), .i2(pp7_w[8 ]), .i3(pp8_w[6 ]), .ci(stg1_co2[11]), .s(stg1_s2[12]), .c(stg1_c2[12]), .co(stg1_co2[12]));
counter_5to3 u_a12_13(.i0(pp5_w[13]), .i1(pp6_w[11]), .i2(pp7_w[9 ]), .i3(pp8_w[7 ]), .ci(stg1_co2[12]), .s(stg1_s2[13]), .c(stg1_c2[13]), .co(stg1_co2[13]));
counter_5to3 u_a12_14(.i0(pp5_w[14]), .i1(pp6_w[12]), .i2(pp7_w[10]), .i3(pp8_w[8 ]), .ci(stg1_co2[13]), .s(stg1_s2[14]), .c(stg1_c2[14]), .co(stg1_co2[14]));
counter_5to3 u_a12_15(.i0(pp5_w[15]), .i1(pp6_w[13]), .i2(pp7_w[11]), .i3(pp8_w[9 ]), .ci(stg1_co2[14]), .s(stg1_s2[15]), .c(stg1_c2[15]), .co(stg1_co2[15]));
counter_5to3 u_a12_16(.i0(pp5_w[16]), .i1(pp6_w[14]), .i2(pp7_w[12]), .i3(pp8_w[10]), .ci(stg1_co2[15]), .s(stg1_s2[16]), .c(stg1_c2[16]), .co(stg1_co2[16]));
counter_5to3 u_a12_17(.i0(pp5_w[17]), .i1(pp6_w[15]), .i2(pp7_w[13]), .i3(pp8_w[11]), .ci(stg1_co2[16]), .s(stg1_s2[17]), .c(stg1_c2[17]), .co(stg1_co2[17]));
counter_5to3 u_a12_18(.i0(pp5_w[18]), .i1(pp6_w[16]), .i2(pp7_w[14]), .i3(pp8_w[12]), .ci(stg1_co2[17]), .s(stg1_s2[18]), .c(stg1_c2[18]), .co(stg1_co2[18]));
counter_5to3 u_a12_19(.i0(pp5_w[19]), .i1(pp6_w[17]), .i2(pp7_w[15]), .i3(pp8_w[13]), .ci(stg1_co2[18]), .s(stg1_s2[19]), .c(stg1_c2[19]), .co(stg1_co2[19]));
counter_5to3 u_a12_20(.i0(pp5_w[20]), .i1(pp6_w[18]), .i2(pp7_w[16]), .i3(pp8_w[14]), .ci(stg1_co2[19]), .s(stg1_s2[20]), .c(stg1_c2[20]), .co(stg1_co2[20]));
counter_5to3 u_a12_21(.i0(pp5_w[21]), .i1(pp6_w[19]), .i2(pp7_w[17]), .i3(pp8_w[15]), .ci(stg1_co2[20]), .s(stg1_s2[21]), .c(stg1_c2[21]), .co(stg1_co2[21]));
counter_5to3 u_a12_22(.i0(pp5_w[22]), .i1(pp6_w[20]), .i2(pp7_w[18]), .i3(pp8_w[16]), .ci(stg1_co2[21]), .s(stg1_s2[22]), .c(stg1_c2[22]), .co(stg1_co2[22]));
counter_5to3 u_a12_23(.i0(pp5_w[23]), .i1(pp6_w[21]), .i2(pp7_w[19]), .i3(pp8_w[17]), .ci(stg1_co2[22]), .s(stg1_s2[23]), .c(stg1_c2[23]), .co(stg1_co2[23]));
counter_5to3 u_a12_24(.i0(pp5_w[24]), .i1(pp6_w[22]), .i2(pp7_w[20]), .i3(pp8_w[18]), .ci(stg1_co2[23]), .s(stg1_s2[24]), .c(stg1_c2[24]), .co(stg1_co2[24]));
counter_5to3 u_a12_25(.i0(pp5_w[25]), .i1(pp6_w[23]), .i2(pp7_w[21]), .i3(pp8_w[19]), .ci(stg1_co2[24]), .s(stg1_s2[25]), .c(stg1_c2[25]), .co(stg1_co2[25]));
counter_5to3 u_a12_26(.i0(pp5_w[26]), .i1(pp6_w[24]), .i2(pp7_w[22]), .i3(pp8_w[20]), .ci(stg1_co2[25]), .s(stg1_s2[26]), .c(stg1_c2[26]), .co(stg1_co2[26]));
counter_5to3 u_a12_27(.i0(pp5_w[27]), .i1(pp6_w[25]), .i2(pp7_w[23]), .i3(pp8_w[21]), .ci(stg1_co2[26]), .s(stg1_s2[27]), .c(stg1_c2[27]), .co(stg1_co2[27]));
counter_5to3 u_a12_28(.i0(pp5_w[28]), .i1(pp6_w[26]), .i2(pp7_w[24]), .i3(pp8_w[22]), .ci(stg1_co2[27]), .s(stg1_s2[28]), .c(stg1_c2[28]), .co(stg1_co2[28]));
counter_5to3 u_a12_29(.i0(pp5_w[29]), .i1(pp6_w[27]), .i2(pp7_w[25]), .i3(pp8_w[23]), .ci(stg1_co2[28]), .s(stg1_s2[29]), .c(stg1_c2[29]), .co(stg1_co2[29]));
counter_5to3 u_a12_30(.i0(pp5_w[30]), .i1(pp6_w[28]), .i2(pp7_w[26]), .i3(pp8_w[24]), .ci(stg1_co2[29]), .s(stg1_s2[30]), .c(stg1_c2[30]), .co(stg1_co2[30]));
counter_5to3 u_a12_31(.i0(pp5_w[31]), .i1(pp6_w[29]), .i2(pp7_w[27]), .i3(pp8_w[25]), .ci(stg1_co2[30]), .s(stg1_s2[31]), .c(stg1_c2[31]), .co(stg1_co2[31]));
counter_5to3 u_a12_32(.i0(pp5_w[32]), .i1(pp6_w[30]), .i2(pp7_w[28]), .i3(pp8_w[26]), .ci(stg1_co2[31]), .s(stg1_s2[32]), .c(stg1_c2[32]), .co(stg1_co2[32]));
counter_5to3 u_a12_33(.i0(pp5_w[33]), .i1(pp6_w[31]), .i2(pp7_w[29]), .i3(pp8_w[27]), .ci(stg1_co2[32]), .s(stg1_s2[33]), .c(stg1_c2[33]), .co(stg1_co2[33]));
counter_5to3 u_a12_34(.i0(pp5_w[34]), .i1(pp6_w[32]), .i2(pp7_w[30]), .i3(pp8_w[28]), .ci(stg1_co2[33]), .s(stg1_s2[34]), .c(stg1_c2[34]), .co(stg1_co2[34]));
counter_5to3 u_a12_35(.i0(pp5_w[35]), .i1(pp6_w[33]), .i2(pp7_w[31]), .i3(pp8_w[29]), .ci(stg1_co2[34]), .s(stg1_s2[35]), .c(stg1_c2[35]), .co(stg1_co2[35]));
counter_5to3 u_a12_36(.i0(pp5_w[36]), .i1(pp6_w[34]), .i2(pp7_w[32]), .i3(pp8_w[30]), .ci(stg1_co2[35]), .s(stg1_s2[36]), .c(stg1_c2[36]), .co(stg1_co2[36]));
counter_5to3 u_a12_37(.i0(pp5_w[37]), .i1(pp6_w[35]), .i2(pp7_w[33]), .i3(pp8_w[31]), .ci(stg1_co2[36]), .s(stg1_s2[37]), .c(stg1_c2[37]), .co(stg1_co2[37]));
counter_5to3 u_a12_38(.i0(pp5_w[38]), .i1(pp6_w[36]), .i2(pp7_w[34]), .i3(pp8_w[32]), .ci(stg1_co2[37]), .s(stg1_s2[38]), .c(stg1_c2[38]), .co(stg1_co2[38]));
counter_5to3 u_a12_39(.i0(pp5_w[39]), .i1(pp6_w[37]), .i2(pp7_w[35]), .i3(pp8_w[33]), .ci(stg1_co2[38]), .s(stg1_s2[39]), .c(stg1_c2[39]), .co(stg1_co2[39]));
counter_5to3 u_a12_40(.i0(pp5_w[40]), .i1(pp6_w[38]), .i2(pp7_w[36]), .i3(pp8_w[34]), .ci(stg1_co2[39]), .s(stg1_s2[40]), .c(stg1_c2[40]), .co(stg1_co2[40]));
counter_5to3 u_a12_41(.i0(pp5_w[41]), .i1(pp6_w[39]), .i2(pp7_w[37]), .i3(pp8_w[35]), .ci(stg1_co2[40]), .s(stg1_s2[41]), .c(stg1_c2[41]), .co(stg1_co2[41]));
counter_5to3 u_a12_42(.i0(pp5_w[42]), .i1(pp6_w[40]), .i2(pp7_w[38]), .i3(pp8_w[36]), .ci(stg1_co2[41]), .s(stg1_s2[42]), .c(stg1_c2[42]), .co(stg1_co2[42]));
counter_5to3 u_a12_43(.i0(pp5_w[43]), .i1(pp6_w[41]), .i2(pp7_w[39]), .i3(pp8_w[37]), .ci(stg1_co2[42]), .s(stg1_s2[43]), .c(stg1_c2[43]), .co(stg1_co2[43]));
counter_5to3 u_a12_44(.i0(pp5_w[44]), .i1(pp6_w[42]), .i2(pp7_w[40]), .i3(pp8_w[38]), .ci(stg1_co2[43]), .s(stg1_s2[44]), .c(stg1_c2[44]), .co(stg1_co2[44]));
counter_5to3 u_a12_45(.i0(pp5_w[45]), .i1(pp6_w[43]), .i2(pp7_w[41]), .i3(pp8_w[39]), .ci(stg1_co2[44]), .s(stg1_s2[45]), .c(stg1_c2[45]), .co(stg1_co2[45]));
counter_5to3 u_a12_46(.i0(pp5_w[46]), .i1(pp6_w[44]), .i2(pp7_w[42]), .i3(pp8_w[40]), .ci(stg1_co2[45]), .s(stg1_s2[46]), .c(stg1_c2[46]), .co(stg1_co2[46]));
counter_5to3 u_a12_47(.i0(pp5_w[47]), .i1(pp6_w[45]), .i2(pp7_w[43]), .i3(pp8_w[41]), .ci(stg1_co2[46]), .s(stg1_s2[47]), .c(stg1_c2[47]), .co(stg1_co2[47]));
counter_5to3 u_a12_48(.i0(pp5_w[48]), .i1(pp6_w[46]), .i2(pp7_w[44]), .i3(pp8_w[42]), .ci(stg1_co2[47]), .s(stg1_s2[48]), .c(stg1_c2[48]), .co(stg1_co2[48]));
counter_5to3 u_a12_49(.i0(pp5_w[49]), .i1(pp6_w[47]), .i2(pp7_w[45]), .i3(pp8_w[43]), .ci(stg1_co2[48]), .s(stg1_s2[49]), .c(stg1_c2[49]), .co(stg1_co2[49]));
counter_5to3 u_a12_50(.i0(pp5_w[50]), .i1(pp6_w[48]), .i2(pp7_w[46]), .i3(pp8_w[44]), .ci(stg1_co2[49]), .s(stg1_s2[50]), .c(stg1_c2[50]), .co(stg1_co2[50]));
counter_5to3 u_a12_51(.i0(pp5_w[51]), .i1(pp6_w[49]), .i2(pp7_w[47]), .i3(pp8_w[45]), .ci(stg1_co2[50]), .s(stg1_s2[51]), .c(stg1_c2[51]), .co(stg1_co2[51]));
counter_5to3 u_a12_52(.i0(pp5_w[52]), .i1(pp6_w[50]), .i2(pp7_w[48]), .i3(pp8_w[46]), .ci(stg1_co2[51]), .s(stg1_s2[52]), .c(stg1_c2[52]), .co(stg1_co2[52]));
counter_5to3 u_a12_53(.i0(pp5_w[53]), .i1(pp6_w[51]), .i2(pp7_w[49]), .i3(pp8_w[47]), .ci(stg1_co2[52]), .s(stg1_s2[53]), .c(stg1_c2[53]), .co(stg1_co2[53]));
counter_5to3 u_a12_54(.i0(pp5_w[54]), .i1(pp6_w[52]), .i2(pp7_w[50]), .i3(pp8_w[48]), .ci(stg1_co2[53]), .s(stg1_s2[54]), .c(stg1_c2[54]), .co(stg1_co2[54]));
counter_5to3 u_a12_55(.i0(pp5_w[55]), .i1(pp6_w[53]), .i2(pp7_w[51]), .i3(pp8_w[49]), .ci(stg1_co2[54]), .s(stg1_s2[55]), .c(stg1_c2[55]), .co(stg1_co2[55]));
counter_5to3 u_a12_56(.i0(pp5_w[56]), .i1(pp6_w[54]), .i2(pp7_w[52]), .i3(pp8_w[50]), .ci(stg1_co2[55]), .s(stg1_s2[56]), .c(stg1_c2[56]), .co(stg1_co2[56]));
counter_5to3 u_a12_57(.i0(pp5_w[57]), .i1(pp6_w[55]), .i2(pp7_w[53]), .i3(pp8_w[51]), .ci(stg1_co2[56]), .s(stg1_s2[57]), .c(stg1_c2[57]), .co(stg1_co2[57]));
counter_5to3 u_a12_58(.i0(pp5_w[58]), .i1(pp6_w[56]), .i2(pp7_w[54]), .i3(pp8_w[52]), .ci(stg1_co2[57]), .s(stg1_s2[58]), .c(stg1_c2[58]), .co(stg1_co2[58]));
counter_5to3 u_a12_59(.i0(pp5_w[59]), .i1(pp6_w[57]), .i2(pp7_w[55]), .i3(pp8_w[53]), .ci(stg1_co2[58]), .s(stg1_s2[59]), .c(stg1_c2[59]), .co(stg1_co2[59]));
counter_5to3 u_a12_60(.i0(pp5_w[60]), .i1(pp6_w[58]), .i2(pp7_w[56]), .i3(pp8_w[54]), .ci(stg1_co2[59]), .s(stg1_s2[60]), .c(stg1_c2[60]), .co(stg1_co2[60]));
counter_5to3 u_a12_61(.i0(pp5_w[61]), .i1(pp6_w[59]), .i2(pp7_w[57]), .i3(pp8_w[55]), .ci(stg1_co2[60]), .s(stg1_s2[61]), .c(stg1_c2[61]), .co(stg1_co2[61]));
counter_5to3 u_a12_62(.i0(pp5_w[62]), .i1(pp6_w[60]), .i2(pp7_w[58]), .i3(pp8_w[56]), .ci(stg1_co2[61]), .s(stg1_s2[62]), .c(stg1_c2[62]), .co(stg1_co2[62]));
counter_5to3 u_a12_63(.i0(pp5_w[63]), .i1(pp6_w[61]), .i2(pp7_w[59]), .i3(pp8_w[57]), .ci(stg1_co2[62]), .s(stg1_s2[63]), .c(stg1_c2[63]), .co(stg1_co2[63]));
counter_5to3 u_a12_64(.i0(pp5_w[64]), .i1(pp6_w[62]), .i2(pp7_w[60]), .i3(pp8_w[58]), .ci(stg1_co2[63]), .s(stg1_s2[64]), .c(stg1_c2[64]), .co(stg1_co2[64]));
counter_5to3 u_a12_65(.i0(pp5_w[65]), .i1(pp6_w[63]), .i2(pp7_w[61]), .i3(pp8_w[59]), .ci(stg1_co2[64]), .s(stg1_s2[65]), .c(stg1_c2[65]), .co(stg1_co2[65]));
counter_5to3 u_a12_66(.i0(pp5_w[65]), .i1(pp6_w[64]), .i2(pp7_w[62]), .i3(pp8_w[60]), .ci(stg1_co2[65]), .s(stg1_s2[66]), .c(stg1_c2[66]), .co(stg1_co2[66]));
counter_5to3 u_a12_67(.i0(pp5_w[65]), .i1(pp6_w[65]), .i2(pp7_w[63]), .i3(pp8_w[61]), .ci(stg1_co2[66]), .s(stg1_s2[67]), .c(stg1_c2[67]), .co(stg1_co2[67]));
counter_5to3 u_a12_68(.i0(pp5_w[65]), .i1(pp6_w[65]), .i2(pp7_w[64]), .i3(pp8_w[62]), .ci(stg1_co2[67]), .s(stg1_s2[68]), .c(stg1_c2[68]), .co(stg1_co2[68]));
counter_5to3 u_a12_69(.i0(pp5_w[65]), .i1(pp6_w[65]), .i2(pp7_w[65]), .i3(pp8_w[63]), .ci(stg1_co2[68]), .s(stg1_s2[69]), .c(stg1_c2[69]), .co(stg1_co2[69]));
counter_5to3 u_a12_70(.i0(pp5_w[65]), .i1(pp6_w[65]), .i2(pp7_w[65]), .i3(pp8_w[64]), .ci(stg1_co2[69]), .s(stg1_s2[70]), .c(stg1_c2[70]), .co(stg1_co2[70]));
counter_5to3 u_al2_71(.i0(pp5_w[65]), .i1(pp6_w[65]), .i2(pp7_w[65]), .i3(pp8_w[65]), .ci(stg1_co2[70]), .s(stg1_s2[71]), .c(stg1_c2[71]), .co(stg1_co2[71]));
counter_5to3 u_al2_72(.i0(pp5_w[65]), .i1(pp6_w[65]), .i2(pp7_w[65]), .i3(pp8_w[65]), .ci(stg1_co2[71]), .s(stg1_s2[72]), .c(stg1_c2[72]), .co(stg1_co2[72]));

// =========================== first stage 3rd group ============================================================================================================
counter_5to3 u_a13_0 (.i0(pp9_w[0 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(1'b0        ), .s(stg1_s3[0 ]), .c(stg1_c3[0 ]), .co(stg1_co3[0 ]));
counter_5to3 u_a13_1 (.i0(pp9_w[1 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co3[0 ]), .s(stg1_s3[1 ]), .c(stg1_c3[1 ]), .co(stg1_co3[1 ]));
counter_5to3 u_a13_2 (.i0(pp9_w[2 ]), .i1(pp10_w[0 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co3[1 ]), .s(stg1_s3[2 ]), .c(stg1_c3[2 ]), .co(stg1_co3[2 ]));
counter_5to3 u_a13_3 (.i0(pp9_w[3 ]), .i1(pp10_w[1 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co3[2 ]), .s(stg1_s3[3 ]), .c(stg1_c3[3 ]), .co(stg1_co3[3 ]));
counter_5to3 u_a13_4 (.i0(pp9_w[4 ]), .i1(pp10_w[2 ]), .i2(pp11_w[0 ]), .i3(1'b0      ), .ci(stg1_co3[3 ]), .s(stg1_s3[4 ]), .c(stg1_c3[4 ]), .co(stg1_co3[4 ]));
counter_5to3 u_a13_5 (.i0(pp9_w[5 ]), .i1(pp10_w[3 ]), .i2(pp11_w[1 ]), .i3(1'b0      ), .ci(stg1_co3[4 ]), .s(stg1_s3[5 ]), .c(stg1_c3[5 ]), .co(stg1_co3[5 ]));
counter_5to3 u_a13_6 (.i0(pp9_w[6 ]), .i1(pp10_w[4 ]), .i2(pp11_w[2 ]), .i3(pp12_w[0 ]), .ci(stg1_co3[5 ]), .s(stg1_s3[6 ]), .c(stg1_c3[6 ]), .co(stg1_co3[6 ]));
counter_5to3 u_a13_7 (.i0(pp9_w[7 ]), .i1(pp10_w[5 ]), .i2(pp11_w[3 ]), .i3(pp12_w[1 ]), .ci(stg1_co3[6 ]), .s(stg1_s3[7 ]), .c(stg1_c3[7 ]), .co(stg1_co3[7 ]));
counter_5to3 u_a13_8 (.i0(pp9_w[8 ]), .i1(pp10_w[6 ]), .i2(pp11_w[4 ]), .i3(pp12_w[2 ]), .ci(stg1_co3[7 ]), .s(stg1_s3[8 ]), .c(stg1_c3[8 ]), .co(stg1_co3[8 ]));
counter_5to3 u_a13_9 (.i0(pp9_w[9 ]), .i1(pp10_w[7 ]), .i2(pp11_w[5 ]), .i3(pp12_w[3 ]), .ci(stg1_co3[8 ]), .s(stg1_s3[9 ]), .c(stg1_c3[9 ]), .co(stg1_co3[9 ]));
counter_5to3 u_a13_10(.i0(pp9_w[10]), .i1(pp10_w[8 ]), .i2(pp11_w[6 ]), .i3(pp12_w[4 ]), .ci(stg1_co3[9 ]), .s(stg1_s3[10]), .c(stg1_c3[10]), .co(stg1_co3[10]));
counter_5to3 u_a13_11(.i0(pp9_w[11]), .i1(pp10_w[9 ]), .i2(pp11_w[7 ]), .i3(pp12_w[5 ]), .ci(stg1_co3[10]), .s(stg1_s3[11]), .c(stg1_c3[11]), .co(stg1_co3[11]));
counter_5to3 u_a13_12(.i0(pp9_w[12]), .i1(pp10_w[10]), .i2(pp11_w[8 ]), .i3(pp12_w[6 ]), .ci(stg1_co3[11]), .s(stg1_s3[12]), .c(stg1_c3[12]), .co(stg1_co3[12]));
counter_5to3 u_a13_13(.i0(pp9_w[13]), .i1(pp10_w[11]), .i2(pp11_w[9 ]), .i3(pp12_w[7 ]), .ci(stg1_co3[12]), .s(stg1_s3[13]), .c(stg1_c3[13]), .co(stg1_co3[13]));
counter_5to3 u_a13_14(.i0(pp9_w[14]), .i1(pp10_w[12]), .i2(pp11_w[10]), .i3(pp12_w[8 ]), .ci(stg1_co3[13]), .s(stg1_s3[14]), .c(stg1_c3[14]), .co(stg1_co3[14]));
counter_5to3 u_a13_15(.i0(pp9_w[15]), .i1(pp10_w[13]), .i2(pp11_w[11]), .i3(pp12_w[9 ]), .ci(stg1_co3[14]), .s(stg1_s3[15]), .c(stg1_c3[15]), .co(stg1_co3[15]));
counter_5to3 u_a13_16(.i0(pp9_w[16]), .i1(pp10_w[14]), .i2(pp11_w[12]), .i3(pp12_w[10]), .ci(stg1_co3[15]), .s(stg1_s3[16]), .c(stg1_c3[16]), .co(stg1_co3[16]));
counter_5to3 u_a13_17(.i0(pp9_w[17]), .i1(pp10_w[15]), .i2(pp11_w[13]), .i3(pp12_w[11]), .ci(stg1_co3[16]), .s(stg1_s3[17]), .c(stg1_c3[17]), .co(stg1_co3[17]));
counter_5to3 u_a13_18(.i0(pp9_w[18]), .i1(pp10_w[16]), .i2(pp11_w[14]), .i3(pp12_w[12]), .ci(stg1_co3[17]), .s(stg1_s3[18]), .c(stg1_c3[18]), .co(stg1_co3[18]));
counter_5to3 u_a13_19(.i0(pp9_w[19]), .i1(pp10_w[17]), .i2(pp11_w[15]), .i3(pp12_w[13]), .ci(stg1_co3[18]), .s(stg1_s3[19]), .c(stg1_c3[19]), .co(stg1_co3[19]));
counter_5to3 u_a13_20(.i0(pp9_w[20]), .i1(pp10_w[18]), .i2(pp11_w[16]), .i3(pp12_w[14]), .ci(stg1_co3[19]), .s(stg1_s3[20]), .c(stg1_c3[20]), .co(stg1_co3[20]));
counter_5to3 u_a13_21(.i0(pp9_w[21]), .i1(pp10_w[19]), .i2(pp11_w[17]), .i3(pp12_w[15]), .ci(stg1_co3[20]), .s(stg1_s3[21]), .c(stg1_c3[21]), .co(stg1_co3[21]));
counter_5to3 u_a13_22(.i0(pp9_w[22]), .i1(pp10_w[20]), .i2(pp11_w[18]), .i3(pp12_w[16]), .ci(stg1_co3[21]), .s(stg1_s3[22]), .c(stg1_c3[22]), .co(stg1_co3[22]));
counter_5to3 u_a13_23(.i0(pp9_w[23]), .i1(pp10_w[21]), .i2(pp11_w[19]), .i3(pp12_w[17]), .ci(stg1_co3[22]), .s(stg1_s3[23]), .c(stg1_c3[23]), .co(stg1_co3[23]));
counter_5to3 u_a13_24(.i0(pp9_w[24]), .i1(pp10_w[22]), .i2(pp11_w[20]), .i3(pp12_w[18]), .ci(stg1_co3[23]), .s(stg1_s3[24]), .c(stg1_c3[24]), .co(stg1_co3[24]));
counter_5to3 u_a13_25(.i0(pp9_w[25]), .i1(pp10_w[23]), .i2(pp11_w[21]), .i3(pp12_w[19]), .ci(stg1_co3[24]), .s(stg1_s3[25]), .c(stg1_c3[25]), .co(stg1_co3[25]));
counter_5to3 u_a13_26(.i0(pp9_w[26]), .i1(pp10_w[24]), .i2(pp11_w[22]), .i3(pp12_w[20]), .ci(stg1_co3[25]), .s(stg1_s3[26]), .c(stg1_c3[26]), .co(stg1_co3[26]));
counter_5to3 u_a13_27(.i0(pp9_w[27]), .i1(pp10_w[25]), .i2(pp11_w[23]), .i3(pp12_w[21]), .ci(stg1_co3[26]), .s(stg1_s3[27]), .c(stg1_c3[27]), .co(stg1_co3[27]));
counter_5to3 u_a13_28(.i0(pp9_w[28]), .i1(pp10_w[26]), .i2(pp11_w[24]), .i3(pp12_w[22]), .ci(stg1_co3[27]), .s(stg1_s3[28]), .c(stg1_c3[28]), .co(stg1_co3[28]));
counter_5to3 u_a13_29(.i0(pp9_w[29]), .i1(pp10_w[27]), .i2(pp11_w[25]), .i3(pp12_w[23]), .ci(stg1_co3[28]), .s(stg1_s3[29]), .c(stg1_c3[29]), .co(stg1_co3[29]));
counter_5to3 u_a13_30(.i0(pp9_w[30]), .i1(pp10_w[28]), .i2(pp11_w[26]), .i3(pp12_w[24]), .ci(stg1_co3[29]), .s(stg1_s3[30]), .c(stg1_c3[30]), .co(stg1_co3[30]));
counter_5to3 u_a13_31(.i0(pp9_w[31]), .i1(pp10_w[29]), .i2(pp11_w[27]), .i3(pp12_w[25]), .ci(stg1_co3[30]), .s(stg1_s3[31]), .c(stg1_c3[31]), .co(stg1_co3[31]));
counter_5to3 u_a13_32(.i0(pp9_w[32]), .i1(pp10_w[30]), .i2(pp11_w[28]), .i3(pp12_w[26]), .ci(stg1_co3[31]), .s(stg1_s3[32]), .c(stg1_c3[32]), .co(stg1_co3[32]));
counter_5to3 u_a13_33(.i0(pp9_w[33]), .i1(pp10_w[31]), .i2(pp11_w[29]), .i3(pp12_w[27]), .ci(stg1_co3[32]), .s(stg1_s3[33]), .c(stg1_c3[33]), .co(stg1_co3[33]));
counter_5to3 u_a13_34(.i0(pp9_w[34]), .i1(pp10_w[32]), .i2(pp11_w[30]), .i3(pp12_w[28]), .ci(stg1_co3[33]), .s(stg1_s3[34]), .c(stg1_c3[34]), .co(stg1_co3[34]));
counter_5to3 u_a13_35(.i0(pp9_w[35]), .i1(pp10_w[33]), .i2(pp11_w[31]), .i3(pp12_w[29]), .ci(stg1_co3[34]), .s(stg1_s3[35]), .c(stg1_c3[35]), .co(stg1_co3[35]));
counter_5to3 u_a13_36(.i0(pp9_w[36]), .i1(pp10_w[34]), .i2(pp11_w[32]), .i3(pp12_w[30]), .ci(stg1_co3[35]), .s(stg1_s3[36]), .c(stg1_c3[36]), .co(stg1_co3[36]));
counter_5to3 u_a13_37(.i0(pp9_w[37]), .i1(pp10_w[35]), .i2(pp11_w[33]), .i3(pp12_w[31]), .ci(stg1_co3[36]), .s(stg1_s3[37]), .c(stg1_c3[37]), .co(stg1_co3[37]));
counter_5to3 u_a13_38(.i0(pp9_w[38]), .i1(pp10_w[36]), .i2(pp11_w[34]), .i3(pp12_w[32]), .ci(stg1_co3[37]), .s(stg1_s3[38]), .c(stg1_c3[38]), .co(stg1_co3[38]));
counter_5to3 u_a13_39(.i0(pp9_w[39]), .i1(pp10_w[37]), .i2(pp11_w[35]), .i3(pp12_w[33]), .ci(stg1_co3[38]), .s(stg1_s3[39]), .c(stg1_c3[39]), .co(stg1_co3[39]));
counter_5to3 u_a13_40(.i0(pp9_w[40]), .i1(pp10_w[38]), .i2(pp11_w[36]), .i3(pp12_w[34]), .ci(stg1_co3[39]), .s(stg1_s3[40]), .c(stg1_c3[40]), .co(stg1_co3[40]));
counter_5to3 u_a13_41(.i0(pp9_w[41]), .i1(pp10_w[39]), .i2(pp11_w[37]), .i3(pp12_w[35]), .ci(stg1_co3[40]), .s(stg1_s3[41]), .c(stg1_c3[41]), .co(stg1_co3[41]));
counter_5to3 u_a13_42(.i0(pp9_w[42]), .i1(pp10_w[40]), .i2(pp11_w[38]), .i3(pp12_w[36]), .ci(stg1_co3[41]), .s(stg1_s3[42]), .c(stg1_c3[42]), .co(stg1_co3[42]));
counter_5to3 u_a13_43(.i0(pp9_w[43]), .i1(pp10_w[41]), .i2(pp11_w[39]), .i3(pp12_w[37]), .ci(stg1_co3[42]), .s(stg1_s3[43]), .c(stg1_c3[43]), .co(stg1_co3[43]));
counter_5to3 u_a13_44(.i0(pp9_w[44]), .i1(pp10_w[42]), .i2(pp11_w[40]), .i3(pp12_w[38]), .ci(stg1_co3[43]), .s(stg1_s3[44]), .c(stg1_c3[44]), .co(stg1_co3[44]));
counter_5to3 u_a13_45(.i0(pp9_w[45]), .i1(pp10_w[43]), .i2(pp11_w[41]), .i3(pp12_w[39]), .ci(stg1_co3[44]), .s(stg1_s3[45]), .c(stg1_c3[45]), .co(stg1_co3[45]));
counter_5to3 u_a13_46(.i0(pp9_w[46]), .i1(pp10_w[44]), .i2(pp11_w[42]), .i3(pp12_w[40]), .ci(stg1_co3[45]), .s(stg1_s3[46]), .c(stg1_c3[46]), .co(stg1_co3[46]));
counter_5to3 u_a13_47(.i0(pp9_w[47]), .i1(pp10_w[45]), .i2(pp11_w[43]), .i3(pp12_w[41]), .ci(stg1_co3[46]), .s(stg1_s3[47]), .c(stg1_c3[47]), .co(stg1_co3[47]));
counter_5to3 u_a13_48(.i0(pp9_w[48]), .i1(pp10_w[46]), .i2(pp11_w[44]), .i3(pp12_w[42]), .ci(stg1_co3[47]), .s(stg1_s3[48]), .c(stg1_c3[48]), .co(stg1_co3[48]));
counter_5to3 u_a13_49(.i0(pp9_w[49]), .i1(pp10_w[47]), .i2(pp11_w[45]), .i3(pp12_w[43]), .ci(stg1_co3[48]), .s(stg1_s3[49]), .c(stg1_c3[49]), .co(stg1_co3[49]));
counter_5to3 u_a13_50(.i0(pp9_w[50]), .i1(pp10_w[48]), .i2(pp11_w[46]), .i3(pp12_w[44]), .ci(stg1_co3[49]), .s(stg1_s3[50]), .c(stg1_c3[50]), .co(stg1_co3[50]));
counter_5to3 u_a13_51(.i0(pp9_w[51]), .i1(pp10_w[49]), .i2(pp11_w[47]), .i3(pp12_w[45]), .ci(stg1_co3[50]), .s(stg1_s3[51]), .c(stg1_c3[51]), .co(stg1_co3[51]));
counter_5to3 u_a13_52(.i0(pp9_w[52]), .i1(pp10_w[50]), .i2(pp11_w[48]), .i3(pp12_w[46]), .ci(stg1_co3[51]), .s(stg1_s3[52]), .c(stg1_c3[52]), .co(stg1_co3[52]));
counter_5to3 u_a13_53(.i0(pp9_w[53]), .i1(pp10_w[51]), .i2(pp11_w[49]), .i3(pp12_w[47]), .ci(stg1_co3[52]), .s(stg1_s3[53]), .c(stg1_c3[53]), .co(stg1_co3[53]));
counter_5to3 u_a13_54(.i0(pp9_w[54]), .i1(pp10_w[52]), .i2(pp11_w[50]), .i3(pp12_w[48]), .ci(stg1_co3[53]), .s(stg1_s3[54]), .c(stg1_c3[54]), .co(stg1_co3[54]));
counter_5to3 u_a13_55(.i0(pp9_w[55]), .i1(pp10_w[53]), .i2(pp11_w[51]), .i3(pp12_w[49]), .ci(stg1_co3[54]), .s(stg1_s3[55]), .c(stg1_c3[55]), .co(stg1_co3[55]));
counter_5to3 u_a13_56(.i0(pp9_w[56]), .i1(pp10_w[54]), .i2(pp11_w[52]), .i3(pp12_w[50]), .ci(stg1_co3[55]), .s(stg1_s3[56]), .c(stg1_c3[56]), .co(stg1_co3[56]));
counter_5to3 u_a13_57(.i0(pp9_w[57]), .i1(pp10_w[55]), .i2(pp11_w[53]), .i3(pp12_w[51]), .ci(stg1_co3[56]), .s(stg1_s3[57]), .c(stg1_c3[57]), .co(stg1_co3[57]));
counter_5to3 u_a13_58(.i0(pp9_w[58]), .i1(pp10_w[56]), .i2(pp11_w[54]), .i3(pp12_w[52]), .ci(stg1_co3[57]), .s(stg1_s3[58]), .c(stg1_c3[58]), .co(stg1_co3[58]));
counter_5to3 u_a13_59(.i0(pp9_w[59]), .i1(pp10_w[57]), .i2(pp11_w[55]), .i3(pp12_w[53]), .ci(stg1_co3[58]), .s(stg1_s3[59]), .c(stg1_c3[59]), .co(stg1_co3[59]));
counter_5to3 u_a13_60(.i0(pp9_w[60]), .i1(pp10_w[58]), .i2(pp11_w[56]), .i3(pp12_w[54]), .ci(stg1_co3[59]), .s(stg1_s3[60]), .c(stg1_c3[60]), .co(stg1_co3[60]));
counter_5to3 u_a13_61(.i0(pp9_w[61]), .i1(pp10_w[59]), .i2(pp11_w[57]), .i3(pp12_w[55]), .ci(stg1_co3[60]), .s(stg1_s3[61]), .c(stg1_c3[61]), .co(stg1_co3[61]));
counter_5to3 u_a13_62(.i0(pp9_w[62]), .i1(pp10_w[60]), .i2(pp11_w[58]), .i3(pp12_w[56]), .ci(stg1_co3[61]), .s(stg1_s3[62]), .c(stg1_c3[62]), .co(stg1_co3[62]));
counter_5to3 u_a13_63(.i0(pp9_w[63]), .i1(pp10_w[61]), .i2(pp11_w[59]), .i3(pp12_w[57]), .ci(stg1_co3[62]), .s(stg1_s3[63]), .c(stg1_c3[63]), .co(stg1_co3[63]));
counter_5to3 u_a13_64(.i0(pp9_w[64]), .i1(pp10_w[62]), .i2(pp11_w[60]), .i3(pp12_w[58]), .ci(stg1_co3[63]), .s(stg1_s3[64]), .c(stg1_c3[64]), .co(stg1_co3[64]));
counter_5to3 u_a13_65(.i0(pp9_w[65]), .i1(pp10_w[63]), .i2(pp11_w[61]), .i3(pp12_w[59]), .ci(stg1_co3[64]), .s(stg1_s3[65]), .c(stg1_c3[65]), .co(stg1_co3[65]));
counter_5to3 u_a13_66(.i0(pp9_w[65]), .i1(pp10_w[64]), .i2(pp11_w[62]), .i3(pp12_w[60]), .ci(stg1_co3[65]), .s(stg1_s3[66]), .c(stg1_c3[66]), .co(stg1_co3[66]));
counter_5to3 u_a13_67(.i0(pp9_w[65]), .i1(pp10_w[65]), .i2(pp11_w[63]), .i3(pp12_w[61]), .ci(stg1_co3[66]), .s(stg1_s3[67]), .c(stg1_c3[67]), .co(stg1_co3[67]));
counter_5to3 u_a13_68(.i0(pp9_w[65]), .i1(pp10_w[65]), .i2(pp11_w[64]), .i3(pp12_w[62]), .ci(stg1_co3[67]), .s(stg1_s3[68]), .c(stg1_c3[68]), .co(stg1_co3[68]));
counter_5to3 u_a13_69(.i0(pp9_w[65]), .i1(pp10_w[65]), .i2(pp11_w[65]), .i3(pp12_w[63]), .ci(stg1_co3[68]), .s(stg1_s3[69]), .c(stg1_c3[69]), .co(stg1_co3[69]));
counter_5to3 u_a13_70(.i0(pp9_w[65]), .i1(pp10_w[65]), .i2(pp11_w[65]), .i3(pp12_w[64]), .ci(stg1_co3[69]), .s(stg1_s3[70]), .c(stg1_c3[70]), .co(stg1_co3[70]));
counter_5to3 u_al3_71(.i0(pp9_w[65]), .i1(pp10_w[65]), .i2(pp11_w[65]), .i3(pp12_w[65]), .ci(stg1_co3[70]), .s(stg1_s3[71]), .c(stg1_c3[71]), .co(stg1_co3[71]));
counter_5to3 u_al3_72(.i0(pp9_w[65]), .i1(pp10_w[65]), .i2(pp11_w[65]), .i3(pp12_w[65]), .ci(stg1_co3[71]), .s(stg1_s3[72]), .c(stg1_c3[72]), .co(stg1_co3[72]));

// =========================== first stage 4th group ============================================================================================================
counter_5to3 u_a14_0 (.i0(pp13_w[0 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(1'b0        ), .s(stg1_s4[0 ]), .c(stg1_c4[0 ]), .co(stg1_co4[0 ]));
counter_5to3 u_a14_1 (.i0(pp13_w[1 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co4[0 ]), .s(stg1_s4[1 ]), .c(stg1_c4[1 ]), .co(stg1_co4[1 ]));
counter_5to3 u_a14_2 (.i0(pp13_w[2 ]), .i1(pp14_w[0 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co4[1 ]), .s(stg1_s4[2 ]), .c(stg1_c4[2 ]), .co(stg1_co4[2 ]));
counter_5to3 u_a14_3 (.i0(pp13_w[3 ]), .i1(pp14_w[1 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co4[2 ]), .s(stg1_s4[3 ]), .c(stg1_c4[3 ]), .co(stg1_co4[3 ]));
counter_5to3 u_a14_4 (.i0(pp13_w[4 ]), .i1(pp14_w[2 ]), .i2(pp15_w[0 ]), .i3(1'b0      ), .ci(stg1_co4[3 ]), .s(stg1_s4[4 ]), .c(stg1_c4[4 ]), .co(stg1_co4[4 ]));
counter_5to3 u_a14_5 (.i0(pp13_w[5 ]), .i1(pp14_w[3 ]), .i2(pp15_w[1 ]), .i3(1'b0      ), .ci(stg1_co4[4 ]), .s(stg1_s4[5 ]), .c(stg1_c4[5 ]), .co(stg1_co4[5 ]));
counter_5to3 u_a14_6 (.i0(pp13_w[6 ]), .i1(pp14_w[4 ]), .i2(pp15_w[2 ]), .i3(pp16_w[0 ]), .ci(stg1_co4[5 ]), .s(stg1_s4[6 ]), .c(stg1_c4[6 ]), .co(stg1_co4[6 ]));
counter_5to3 u_a14_7 (.i0(pp13_w[7 ]), .i1(pp14_w[5 ]), .i2(pp15_w[3 ]), .i3(pp16_w[1 ]), .ci(stg1_co4[6 ]), .s(stg1_s4[7 ]), .c(stg1_c4[7 ]), .co(stg1_co4[7 ]));
counter_5to3 u_a14_8 (.i0(pp13_w[8 ]), .i1(pp14_w[6 ]), .i2(pp15_w[4 ]), .i3(pp16_w[2 ]), .ci(stg1_co4[7 ]), .s(stg1_s4[8 ]), .c(stg1_c4[8 ]), .co(stg1_co4[8 ]));
counter_5to3 u_a14_9 (.i0(pp13_w[9 ]), .i1(pp14_w[7 ]), .i2(pp15_w[5 ]), .i3(pp16_w[3 ]), .ci(stg1_co4[8 ]), .s(stg1_s4[9 ]), .c(stg1_c4[9 ]), .co(stg1_co4[9 ]));
counter_5to3 u_a14_10(.i0(pp13_w[10]), .i1(pp14_w[8 ]), .i2(pp15_w[6 ]), .i3(pp16_w[4 ]), .ci(stg1_co4[9 ]), .s(stg1_s4[10]), .c(stg1_c4[10]), .co(stg1_co4[10]));
counter_5to3 u_a14_11(.i0(pp13_w[11]), .i1(pp14_w[9 ]), .i2(pp15_w[7 ]), .i3(pp16_w[5 ]), .ci(stg1_co4[10]), .s(stg1_s4[11]), .c(stg1_c4[11]), .co(stg1_co4[11]));
counter_5to3 u_a14_12(.i0(pp13_w[12]), .i1(pp14_w[10]), .i2(pp15_w[8 ]), .i3(pp16_w[6 ]), .ci(stg1_co4[11]), .s(stg1_s4[12]), .c(stg1_c4[12]), .co(stg1_co4[12]));
counter_5to3 u_a14_13(.i0(pp13_w[13]), .i1(pp14_w[11]), .i2(pp15_w[9 ]), .i3(pp16_w[7 ]), .ci(stg1_co4[12]), .s(stg1_s4[13]), .c(stg1_c4[13]), .co(stg1_co4[13]));
counter_5to3 u_a14_14(.i0(pp13_w[14]), .i1(pp14_w[12]), .i2(pp15_w[10]), .i3(pp16_w[8 ]), .ci(stg1_co4[13]), .s(stg1_s4[14]), .c(stg1_c4[14]), .co(stg1_co4[14]));
counter_5to3 u_a14_15(.i0(pp13_w[15]), .i1(pp14_w[13]), .i2(pp15_w[11]), .i3(pp16_w[9 ]), .ci(stg1_co4[14]), .s(stg1_s4[15]), .c(stg1_c4[15]), .co(stg1_co4[15]));
counter_5to3 u_a14_16(.i0(pp13_w[16]), .i1(pp14_w[14]), .i2(pp15_w[12]), .i3(pp16_w[10]), .ci(stg1_co4[15]), .s(stg1_s4[16]), .c(stg1_c4[16]), .co(stg1_co4[16]));
counter_5to3 u_a14_17(.i0(pp13_w[17]), .i1(pp14_w[15]), .i2(pp15_w[13]), .i3(pp16_w[11]), .ci(stg1_co4[16]), .s(stg1_s4[17]), .c(stg1_c4[17]), .co(stg1_co4[17]));
counter_5to3 u_a14_18(.i0(pp13_w[18]), .i1(pp14_w[16]), .i2(pp15_w[14]), .i3(pp16_w[12]), .ci(stg1_co4[17]), .s(stg1_s4[18]), .c(stg1_c4[18]), .co(stg1_co4[18]));
counter_5to3 u_a14_19(.i0(pp13_w[19]), .i1(pp14_w[17]), .i2(pp15_w[15]), .i3(pp16_w[13]), .ci(stg1_co4[18]), .s(stg1_s4[19]), .c(stg1_c4[19]), .co(stg1_co4[19]));
counter_5to3 u_a14_20(.i0(pp13_w[20]), .i1(pp14_w[18]), .i2(pp15_w[16]), .i3(pp16_w[14]), .ci(stg1_co4[19]), .s(stg1_s4[20]), .c(stg1_c4[20]), .co(stg1_co4[20]));
counter_5to3 u_a14_21(.i0(pp13_w[21]), .i1(pp14_w[19]), .i2(pp15_w[17]), .i3(pp16_w[15]), .ci(stg1_co4[20]), .s(stg1_s4[21]), .c(stg1_c4[21]), .co(stg1_co4[21]));
counter_5to3 u_a14_22(.i0(pp13_w[22]), .i1(pp14_w[20]), .i2(pp15_w[18]), .i3(pp16_w[16]), .ci(stg1_co4[21]), .s(stg1_s4[22]), .c(stg1_c4[22]), .co(stg1_co4[22]));
counter_5to3 u_a14_23(.i0(pp13_w[23]), .i1(pp14_w[21]), .i2(pp15_w[19]), .i3(pp16_w[17]), .ci(stg1_co4[22]), .s(stg1_s4[23]), .c(stg1_c4[23]), .co(stg1_co4[23]));
counter_5to3 u_a14_24(.i0(pp13_w[24]), .i1(pp14_w[22]), .i2(pp15_w[20]), .i3(pp16_w[18]), .ci(stg1_co4[23]), .s(stg1_s4[24]), .c(stg1_c4[24]), .co(stg1_co4[24]));
counter_5to3 u_a14_25(.i0(pp13_w[25]), .i1(pp14_w[23]), .i2(pp15_w[21]), .i3(pp16_w[19]), .ci(stg1_co4[24]), .s(stg1_s4[25]), .c(stg1_c4[25]), .co(stg1_co4[25]));
counter_5to3 u_a14_26(.i0(pp13_w[26]), .i1(pp14_w[24]), .i2(pp15_w[22]), .i3(pp16_w[20]), .ci(stg1_co4[25]), .s(stg1_s4[26]), .c(stg1_c4[26]), .co(stg1_co4[26]));
counter_5to3 u_a14_27(.i0(pp13_w[27]), .i1(pp14_w[25]), .i2(pp15_w[23]), .i3(pp16_w[21]), .ci(stg1_co4[26]), .s(stg1_s4[27]), .c(stg1_c4[27]), .co(stg1_co4[27]));
counter_5to3 u_a14_28(.i0(pp13_w[28]), .i1(pp14_w[26]), .i2(pp15_w[24]), .i3(pp16_w[22]), .ci(stg1_co4[27]), .s(stg1_s4[28]), .c(stg1_c4[28]), .co(stg1_co4[28]));
counter_5to3 u_a14_29(.i0(pp13_w[29]), .i1(pp14_w[27]), .i2(pp15_w[25]), .i3(pp16_w[23]), .ci(stg1_co4[28]), .s(stg1_s4[29]), .c(stg1_c4[29]), .co(stg1_co4[29]));
counter_5to3 u_a14_30(.i0(pp13_w[30]), .i1(pp14_w[28]), .i2(pp15_w[26]), .i3(pp16_w[24]), .ci(stg1_co4[29]), .s(stg1_s4[30]), .c(stg1_c4[30]), .co(stg1_co4[30]));
counter_5to3 u_a14_31(.i0(pp13_w[31]), .i1(pp14_w[29]), .i2(pp15_w[27]), .i3(pp16_w[25]), .ci(stg1_co4[30]), .s(stg1_s4[31]), .c(stg1_c4[31]), .co(stg1_co4[31]));
counter_5to3 u_a14_32(.i0(pp13_w[32]), .i1(pp14_w[30]), .i2(pp15_w[28]), .i3(pp16_w[26]), .ci(stg1_co4[31]), .s(stg1_s4[32]), .c(stg1_c4[32]), .co(stg1_co4[32]));
counter_5to3 u_a14_33(.i0(pp13_w[33]), .i1(pp14_w[31]), .i2(pp15_w[29]), .i3(pp16_w[27]), .ci(stg1_co4[32]), .s(stg1_s4[33]), .c(stg1_c4[33]), .co(stg1_co4[33]));
counter_5to3 u_a14_34(.i0(pp13_w[34]), .i1(pp14_w[32]), .i2(pp15_w[30]), .i3(pp16_w[28]), .ci(stg1_co4[33]), .s(stg1_s4[34]), .c(stg1_c4[34]), .co(stg1_co4[34]));
counter_5to3 u_a14_35(.i0(pp13_w[35]), .i1(pp14_w[33]), .i2(pp15_w[31]), .i3(pp16_w[29]), .ci(stg1_co4[34]), .s(stg1_s4[35]), .c(stg1_c4[35]), .co(stg1_co4[35]));
counter_5to3 u_a14_36(.i0(pp13_w[36]), .i1(pp14_w[34]), .i2(pp15_w[32]), .i3(pp16_w[30]), .ci(stg1_co4[35]), .s(stg1_s4[36]), .c(stg1_c4[36]), .co(stg1_co4[36]));
counter_5to3 u_a14_37(.i0(pp13_w[37]), .i1(pp14_w[35]), .i2(pp15_w[33]), .i3(pp16_w[31]), .ci(stg1_co4[36]), .s(stg1_s4[37]), .c(stg1_c4[37]), .co(stg1_co4[37]));
counter_5to3 u_a14_38(.i0(pp13_w[38]), .i1(pp14_w[36]), .i2(pp15_w[34]), .i3(pp16_w[32]), .ci(stg1_co4[37]), .s(stg1_s4[38]), .c(stg1_c4[38]), .co(stg1_co4[38]));
counter_5to3 u_a14_39(.i0(pp13_w[39]), .i1(pp14_w[37]), .i2(pp15_w[35]), .i3(pp16_w[33]), .ci(stg1_co4[38]), .s(stg1_s4[39]), .c(stg1_c4[39]), .co(stg1_co4[39]));
counter_5to3 u_a14_40(.i0(pp13_w[40]), .i1(pp14_w[38]), .i2(pp15_w[36]), .i3(pp16_w[34]), .ci(stg1_co4[39]), .s(stg1_s4[40]), .c(stg1_c4[40]), .co(stg1_co4[40]));
counter_5to3 u_a14_41(.i0(pp13_w[41]), .i1(pp14_w[39]), .i2(pp15_w[37]), .i3(pp16_w[35]), .ci(stg1_co4[40]), .s(stg1_s4[41]), .c(stg1_c4[41]), .co(stg1_co4[41]));
counter_5to3 u_a14_42(.i0(pp13_w[42]), .i1(pp14_w[40]), .i2(pp15_w[38]), .i3(pp16_w[36]), .ci(stg1_co4[41]), .s(stg1_s4[42]), .c(stg1_c4[42]), .co(stg1_co4[42]));
counter_5to3 u_a14_43(.i0(pp13_w[43]), .i1(pp14_w[41]), .i2(pp15_w[39]), .i3(pp16_w[37]), .ci(stg1_co4[42]), .s(stg1_s4[43]), .c(stg1_c4[43]), .co(stg1_co4[43]));
counter_5to3 u_a14_44(.i0(pp13_w[44]), .i1(pp14_w[42]), .i2(pp15_w[40]), .i3(pp16_w[38]), .ci(stg1_co4[43]), .s(stg1_s4[44]), .c(stg1_c4[44]), .co(stg1_co4[44]));
counter_5to3 u_a14_45(.i0(pp13_w[45]), .i1(pp14_w[43]), .i2(pp15_w[41]), .i3(pp16_w[39]), .ci(stg1_co4[44]), .s(stg1_s4[45]), .c(stg1_c4[45]), .co(stg1_co4[45]));
counter_5to3 u_a14_46(.i0(pp13_w[46]), .i1(pp14_w[44]), .i2(pp15_w[42]), .i3(pp16_w[40]), .ci(stg1_co4[45]), .s(stg1_s4[46]), .c(stg1_c4[46]), .co(stg1_co4[46]));
counter_5to3 u_a14_47(.i0(pp13_w[47]), .i1(pp14_w[45]), .i2(pp15_w[43]), .i3(pp16_w[41]), .ci(stg1_co4[46]), .s(stg1_s4[47]), .c(stg1_c4[47]), .co(stg1_co4[47]));
counter_5to3 u_a14_48(.i0(pp13_w[48]), .i1(pp14_w[46]), .i2(pp15_w[44]), .i3(pp16_w[42]), .ci(stg1_co4[47]), .s(stg1_s4[48]), .c(stg1_c4[48]), .co(stg1_co4[48]));
counter_5to3 u_a14_49(.i0(pp13_w[49]), .i1(pp14_w[47]), .i2(pp15_w[45]), .i3(pp16_w[43]), .ci(stg1_co4[48]), .s(stg1_s4[49]), .c(stg1_c4[49]), .co(stg1_co4[49]));
counter_5to3 u_a14_50(.i0(pp13_w[50]), .i1(pp14_w[48]), .i2(pp15_w[46]), .i3(pp16_w[44]), .ci(stg1_co4[49]), .s(stg1_s4[50]), .c(stg1_c4[50]), .co(stg1_co4[50]));
counter_5to3 u_a14_51(.i0(pp13_w[51]), .i1(pp14_w[49]), .i2(pp15_w[47]), .i3(pp16_w[45]), .ci(stg1_co4[50]), .s(stg1_s4[51]), .c(stg1_c4[51]), .co(stg1_co4[51]));
counter_5to3 u_a14_52(.i0(pp13_w[52]), .i1(pp14_w[50]), .i2(pp15_w[48]), .i3(pp16_w[46]), .ci(stg1_co4[51]), .s(stg1_s4[52]), .c(stg1_c4[52]), .co(stg1_co4[52]));
counter_5to3 u_a14_53(.i0(pp13_w[53]), .i1(pp14_w[51]), .i2(pp15_w[49]), .i3(pp16_w[47]), .ci(stg1_co4[52]), .s(stg1_s4[53]), .c(stg1_c4[53]), .co(stg1_co4[53]));
counter_5to3 u_a14_54(.i0(pp13_w[54]), .i1(pp14_w[52]), .i2(pp15_w[50]), .i3(pp16_w[48]), .ci(stg1_co4[53]), .s(stg1_s4[54]), .c(stg1_c4[54]), .co(stg1_co4[54]));
counter_5to3 u_a14_55(.i0(pp13_w[55]), .i1(pp14_w[53]), .i2(pp15_w[51]), .i3(pp16_w[49]), .ci(stg1_co4[54]), .s(stg1_s4[55]), .c(stg1_c4[55]), .co(stg1_co4[55]));
counter_5to3 u_a14_56(.i0(pp13_w[56]), .i1(pp14_w[54]), .i2(pp15_w[52]), .i3(pp16_w[50]), .ci(stg1_co4[55]), .s(stg1_s4[56]), .c(stg1_c4[56]), .co(stg1_co4[56]));
counter_5to3 u_a14_57(.i0(pp13_w[57]), .i1(pp14_w[55]), .i2(pp15_w[53]), .i3(pp16_w[51]), .ci(stg1_co4[56]), .s(stg1_s4[57]), .c(stg1_c4[57]), .co(stg1_co4[57]));
counter_5to3 u_a14_58(.i0(pp13_w[58]), .i1(pp14_w[56]), .i2(pp15_w[54]), .i3(pp16_w[52]), .ci(stg1_co4[57]), .s(stg1_s4[58]), .c(stg1_c4[58]), .co(stg1_co4[58]));
counter_5to3 u_a14_59(.i0(pp13_w[59]), .i1(pp14_w[57]), .i2(pp15_w[55]), .i3(pp16_w[53]), .ci(stg1_co4[58]), .s(stg1_s4[59]), .c(stg1_c4[59]), .co(stg1_co4[59]));
counter_5to3 u_a14_60(.i0(pp13_w[60]), .i1(pp14_w[58]), .i2(pp15_w[56]), .i3(pp16_w[54]), .ci(stg1_co4[59]), .s(stg1_s4[60]), .c(stg1_c4[60]), .co(stg1_co4[60]));
counter_5to3 u_a14_61(.i0(pp13_w[61]), .i1(pp14_w[59]), .i2(pp15_w[57]), .i3(pp16_w[55]), .ci(stg1_co4[60]), .s(stg1_s4[61]), .c(stg1_c4[61]), .co(stg1_co4[61]));
counter_5to3 u_a14_62(.i0(pp13_w[62]), .i1(pp14_w[60]), .i2(pp15_w[58]), .i3(pp16_w[56]), .ci(stg1_co4[61]), .s(stg1_s4[62]), .c(stg1_c4[62]), .co(stg1_co4[62]));
counter_5to3 u_a14_63(.i0(pp13_w[63]), .i1(pp14_w[61]), .i2(pp15_w[59]), .i3(pp16_w[57]), .ci(stg1_co4[62]), .s(stg1_s4[63]), .c(stg1_c4[63]), .co(stg1_co4[63]));
counter_5to3 u_a14_64(.i0(pp13_w[64]), .i1(pp14_w[62]), .i2(pp15_w[60]), .i3(pp16_w[58]), .ci(stg1_co4[63]), .s(stg1_s4[64]), .c(stg1_c4[64]), .co(stg1_co4[64]));
counter_5to3 u_a14_65(.i0(pp13_w[65]), .i1(pp14_w[63]), .i2(pp15_w[61]), .i3(pp16_w[59]), .ci(stg1_co4[64]), .s(stg1_s4[65]), .c(stg1_c4[65]), .co(stg1_co4[65]));
counter_5to3 u_a14_66(.i0(pp13_w[65]), .i1(pp14_w[64]), .i2(pp15_w[62]), .i3(pp16_w[60]), .ci(stg1_co4[65]), .s(stg1_s4[66]), .c(stg1_c4[66]), .co(stg1_co4[66]));
counter_5to3 u_a14_67(.i0(pp13_w[65]), .i1(pp14_w[65]), .i2(pp15_w[63]), .i3(pp16_w[61]), .ci(stg1_co4[66]), .s(stg1_s4[67]), .c(stg1_c4[67]), .co(stg1_co4[67]));
counter_5to3 u_a14_68(.i0(pp13_w[65]), .i1(pp14_w[65]), .i2(pp15_w[64]), .i3(pp16_w[62]), .ci(stg1_co4[67]), .s(stg1_s4[68]), .c(stg1_c4[68]), .co(stg1_co4[68]));
counter_5to3 u_a14_69(.i0(pp13_w[65]), .i1(pp14_w[65]), .i2(pp15_w[65]), .i3(pp16_w[63]), .ci(stg1_co4[68]), .s(stg1_s4[69]), .c(stg1_c4[69]), .co(stg1_co4[69]));
counter_5to3 u_a14_70(.i0(pp13_w[65]), .i1(pp14_w[65]), .i2(pp15_w[65]), .i3(pp16_w[64]), .ci(stg1_co4[69]), .s(stg1_s4[70]), .c(stg1_c4[70]), .co(stg1_co4[70]));
counter_5to3 u_al4_71(.i0(pp13_w[65]), .i1(pp14_w[65]), .i2(pp15_w[65]), .i3(pp16_w[65]), .ci(stg1_co4[70]), .s(stg1_s4[71]), .c(stg1_c4[71]), .co(stg1_co4[71]));
counter_5to3 u_al4_72(.i0(pp13_w[65]), .i1(pp14_w[65]), .i2(pp15_w[65]), .i3(pp16_w[65]), .ci(stg1_co4[71]), .s(stg1_s4[72]), .c(stg1_c4[72]), .co(stg1_co4[72]));

// =========================== first stage 5th group ============================================================================================================
counter_5to3 u_a15_0 (.i0(pp17_w[0 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(1'b0        ), .s(stg1_s5[0 ]), .c(stg1_c5[0 ]), .co(stg1_co5[0 ]));
counter_5to3 u_a15_1 (.i0(pp17_w[1 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co5[0 ]), .s(stg1_s5[1 ]), .c(stg1_c5[1 ]), .co(stg1_co5[1 ]));
counter_5to3 u_a15_2 (.i0(pp17_w[2 ]), .i1(pp18_w[0 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co5[1 ]), .s(stg1_s5[2 ]), .c(stg1_c5[2 ]), .co(stg1_co5[2 ]));
counter_5to3 u_a15_3 (.i0(pp17_w[3 ]), .i1(pp18_w[1 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co5[2 ]), .s(stg1_s5[3 ]), .c(stg1_c5[3 ]), .co(stg1_co5[3 ]));
counter_5to3 u_a15_4 (.i0(pp17_w[4 ]), .i1(pp18_w[2 ]), .i2(pp19_w[0 ]), .i3(1'b0      ), .ci(stg1_co5[3 ]), .s(stg1_s5[4 ]), .c(stg1_c5[4 ]), .co(stg1_co5[4 ]));
counter_5to3 u_a15_5 (.i0(pp17_w[5 ]), .i1(pp18_w[3 ]), .i2(pp19_w[1 ]), .i3(1'b0      ), .ci(stg1_co5[4 ]), .s(stg1_s5[5 ]), .c(stg1_c5[5 ]), .co(stg1_co5[5 ]));
counter_5to3 u_a15_6 (.i0(pp17_w[6 ]), .i1(pp18_w[4 ]), .i2(pp19_w[2 ]), .i3(pp20_w[0 ]), .ci(stg1_co5[5 ]), .s(stg1_s5[6 ]), .c(stg1_c5[6 ]), .co(stg1_co5[6 ]));
counter_5to3 u_a15_7 (.i0(pp17_w[7 ]), .i1(pp18_w[5 ]), .i2(pp19_w[3 ]), .i3(pp20_w[1 ]), .ci(stg1_co5[6 ]), .s(stg1_s5[7 ]), .c(stg1_c5[7 ]), .co(stg1_co5[7 ]));
counter_5to3 u_a15_8 (.i0(pp17_w[8 ]), .i1(pp18_w[6 ]), .i2(pp19_w[4 ]), .i3(pp20_w[2 ]), .ci(stg1_co5[7 ]), .s(stg1_s5[8 ]), .c(stg1_c5[8 ]), .co(stg1_co5[8 ]));
counter_5to3 u_a15_9 (.i0(pp17_w[9 ]), .i1(pp18_w[7 ]), .i2(pp19_w[5 ]), .i3(pp20_w[3 ]), .ci(stg1_co5[8 ]), .s(stg1_s5[9 ]), .c(stg1_c5[9 ]), .co(stg1_co5[9 ]));
counter_5to3 u_a15_10(.i0(pp17_w[10]), .i1(pp18_w[8 ]), .i2(pp19_w[6 ]), .i3(pp20_w[4 ]), .ci(stg1_co5[9 ]), .s(stg1_s5[10]), .c(stg1_c5[10]), .co(stg1_co5[10]));
counter_5to3 u_a15_11(.i0(pp17_w[11]), .i1(pp18_w[9 ]), .i2(pp19_w[7 ]), .i3(pp20_w[5 ]), .ci(stg1_co5[10]), .s(stg1_s5[11]), .c(stg1_c5[11]), .co(stg1_co5[11]));
counter_5to3 u_a15_12(.i0(pp17_w[12]), .i1(pp18_w[10]), .i2(pp19_w[8 ]), .i3(pp20_w[6 ]), .ci(stg1_co5[11]), .s(stg1_s5[12]), .c(stg1_c5[12]), .co(stg1_co5[12]));
counter_5to3 u_a15_13(.i0(pp17_w[13]), .i1(pp18_w[11]), .i2(pp19_w[9 ]), .i3(pp20_w[7 ]), .ci(stg1_co5[12]), .s(stg1_s5[13]), .c(stg1_c5[13]), .co(stg1_co5[13]));
counter_5to3 u_a15_14(.i0(pp17_w[14]), .i1(pp18_w[12]), .i2(pp19_w[10]), .i3(pp20_w[8 ]), .ci(stg1_co5[13]), .s(stg1_s5[14]), .c(stg1_c5[14]), .co(stg1_co5[14]));
counter_5to3 u_a15_15(.i0(pp17_w[15]), .i1(pp18_w[13]), .i2(pp19_w[11]), .i3(pp20_w[9 ]), .ci(stg1_co5[14]), .s(stg1_s5[15]), .c(stg1_c5[15]), .co(stg1_co5[15]));
counter_5to3 u_a15_16(.i0(pp17_w[16]), .i1(pp18_w[14]), .i2(pp19_w[12]), .i3(pp20_w[10]), .ci(stg1_co5[15]), .s(stg1_s5[16]), .c(stg1_c5[16]), .co(stg1_co5[16]));
counter_5to3 u_a15_17(.i0(pp17_w[17]), .i1(pp18_w[15]), .i2(pp19_w[13]), .i3(pp20_w[11]), .ci(stg1_co5[16]), .s(stg1_s5[17]), .c(stg1_c5[17]), .co(stg1_co5[17]));
counter_5to3 u_a15_18(.i0(pp17_w[18]), .i1(pp18_w[16]), .i2(pp19_w[14]), .i3(pp20_w[12]), .ci(stg1_co5[17]), .s(stg1_s5[18]), .c(stg1_c5[18]), .co(stg1_co5[18]));
counter_5to3 u_a15_19(.i0(pp17_w[19]), .i1(pp18_w[17]), .i2(pp19_w[15]), .i3(pp20_w[13]), .ci(stg1_co5[18]), .s(stg1_s5[19]), .c(stg1_c5[19]), .co(stg1_co5[19]));
counter_5to3 u_a15_20(.i0(pp17_w[20]), .i1(pp18_w[18]), .i2(pp19_w[16]), .i3(pp20_w[14]), .ci(stg1_co5[19]), .s(stg1_s5[20]), .c(stg1_c5[20]), .co(stg1_co5[20]));
counter_5to3 u_a15_21(.i0(pp17_w[21]), .i1(pp18_w[19]), .i2(pp19_w[17]), .i3(pp20_w[15]), .ci(stg1_co5[20]), .s(stg1_s5[21]), .c(stg1_c5[21]), .co(stg1_co5[21]));
counter_5to3 u_a15_22(.i0(pp17_w[22]), .i1(pp18_w[20]), .i2(pp19_w[18]), .i3(pp20_w[16]), .ci(stg1_co5[21]), .s(stg1_s5[22]), .c(stg1_c5[22]), .co(stg1_co5[22]));
counter_5to3 u_a15_23(.i0(pp17_w[23]), .i1(pp18_w[21]), .i2(pp19_w[19]), .i3(pp20_w[17]), .ci(stg1_co5[22]), .s(stg1_s5[23]), .c(stg1_c5[23]), .co(stg1_co5[23]));
counter_5to3 u_a15_24(.i0(pp17_w[24]), .i1(pp18_w[22]), .i2(pp19_w[20]), .i3(pp20_w[18]), .ci(stg1_co5[23]), .s(stg1_s5[24]), .c(stg1_c5[24]), .co(stg1_co5[24]));
counter_5to3 u_a15_25(.i0(pp17_w[25]), .i1(pp18_w[23]), .i2(pp19_w[21]), .i3(pp20_w[19]), .ci(stg1_co5[24]), .s(stg1_s5[25]), .c(stg1_c5[25]), .co(stg1_co5[25]));
counter_5to3 u_a15_26(.i0(pp17_w[26]), .i1(pp18_w[24]), .i2(pp19_w[22]), .i3(pp20_w[20]), .ci(stg1_co5[25]), .s(stg1_s5[26]), .c(stg1_c5[26]), .co(stg1_co5[26]));
counter_5to3 u_a15_27(.i0(pp17_w[27]), .i1(pp18_w[25]), .i2(pp19_w[23]), .i3(pp20_w[21]), .ci(stg1_co5[26]), .s(stg1_s5[27]), .c(stg1_c5[27]), .co(stg1_co5[27]));
counter_5to3 u_a15_28(.i0(pp17_w[28]), .i1(pp18_w[26]), .i2(pp19_w[24]), .i3(pp20_w[22]), .ci(stg1_co5[27]), .s(stg1_s5[28]), .c(stg1_c5[28]), .co(stg1_co5[28]));
counter_5to3 u_a15_29(.i0(pp17_w[29]), .i1(pp18_w[27]), .i2(pp19_w[25]), .i3(pp20_w[23]), .ci(stg1_co5[28]), .s(stg1_s5[29]), .c(stg1_c5[29]), .co(stg1_co5[29]));
counter_5to3 u_a15_30(.i0(pp17_w[30]), .i1(pp18_w[28]), .i2(pp19_w[26]), .i3(pp20_w[24]), .ci(stg1_co5[29]), .s(stg1_s5[30]), .c(stg1_c5[30]), .co(stg1_co5[30]));
counter_5to3 u_a15_31(.i0(pp17_w[31]), .i1(pp18_w[29]), .i2(pp19_w[27]), .i3(pp20_w[25]), .ci(stg1_co5[30]), .s(stg1_s5[31]), .c(stg1_c5[31]), .co(stg1_co5[31]));
counter_5to3 u_a15_32(.i0(pp17_w[32]), .i1(pp18_w[30]), .i2(pp19_w[28]), .i3(pp20_w[26]), .ci(stg1_co5[31]), .s(stg1_s5[32]), .c(stg1_c5[32]), .co(stg1_co5[32]));
counter_5to3 u_a15_33(.i0(pp17_w[33]), .i1(pp18_w[31]), .i2(pp19_w[29]), .i3(pp20_w[27]), .ci(stg1_co5[32]), .s(stg1_s5[33]), .c(stg1_c5[33]), .co(stg1_co5[33]));
counter_5to3 u_a15_34(.i0(pp17_w[34]), .i1(pp18_w[32]), .i2(pp19_w[30]), .i3(pp20_w[28]), .ci(stg1_co5[33]), .s(stg1_s5[34]), .c(stg1_c5[34]), .co(stg1_co5[34]));
counter_5to3 u_a15_35(.i0(pp17_w[35]), .i1(pp18_w[33]), .i2(pp19_w[31]), .i3(pp20_w[29]), .ci(stg1_co5[34]), .s(stg1_s5[35]), .c(stg1_c5[35]), .co(stg1_co5[35]));
counter_5to3 u_a15_36(.i0(pp17_w[36]), .i1(pp18_w[34]), .i2(pp19_w[32]), .i3(pp20_w[30]), .ci(stg1_co5[35]), .s(stg1_s5[36]), .c(stg1_c5[36]), .co(stg1_co5[36]));
counter_5to3 u_a15_37(.i0(pp17_w[37]), .i1(pp18_w[35]), .i2(pp19_w[33]), .i3(pp20_w[31]), .ci(stg1_co5[36]), .s(stg1_s5[37]), .c(stg1_c5[37]), .co(stg1_co5[37]));
counter_5to3 u_a15_38(.i0(pp17_w[38]), .i1(pp18_w[36]), .i2(pp19_w[34]), .i3(pp20_w[32]), .ci(stg1_co5[37]), .s(stg1_s5[38]), .c(stg1_c5[38]), .co(stg1_co5[38]));
counter_5to3 u_a15_39(.i0(pp17_w[39]), .i1(pp18_w[37]), .i2(pp19_w[35]), .i3(pp20_w[33]), .ci(stg1_co5[38]), .s(stg1_s5[39]), .c(stg1_c5[39]), .co(stg1_co5[39]));
counter_5to3 u_a15_40(.i0(pp17_w[40]), .i1(pp18_w[38]), .i2(pp19_w[36]), .i3(pp20_w[34]), .ci(stg1_co5[39]), .s(stg1_s5[40]), .c(stg1_c5[40]), .co(stg1_co5[40]));
counter_5to3 u_a15_41(.i0(pp17_w[41]), .i1(pp18_w[39]), .i2(pp19_w[37]), .i3(pp20_w[35]), .ci(stg1_co5[40]), .s(stg1_s5[41]), .c(stg1_c5[41]), .co(stg1_co5[41]));
counter_5to3 u_a15_42(.i0(pp17_w[42]), .i1(pp18_w[40]), .i2(pp19_w[38]), .i3(pp20_w[36]), .ci(stg1_co5[41]), .s(stg1_s5[42]), .c(stg1_c5[42]), .co(stg1_co5[42]));
counter_5to3 u_a15_43(.i0(pp17_w[43]), .i1(pp18_w[41]), .i2(pp19_w[39]), .i3(pp20_w[37]), .ci(stg1_co5[42]), .s(stg1_s5[43]), .c(stg1_c5[43]), .co(stg1_co5[43]));
counter_5to3 u_a15_44(.i0(pp17_w[44]), .i1(pp18_w[42]), .i2(pp19_w[40]), .i3(pp20_w[38]), .ci(stg1_co5[43]), .s(stg1_s5[44]), .c(stg1_c5[44]), .co(stg1_co5[44]));
counter_5to3 u_a15_45(.i0(pp17_w[45]), .i1(pp18_w[43]), .i2(pp19_w[41]), .i3(pp20_w[39]), .ci(stg1_co5[44]), .s(stg1_s5[45]), .c(stg1_c5[45]), .co(stg1_co5[45]));
counter_5to3 u_a15_46(.i0(pp17_w[46]), .i1(pp18_w[44]), .i2(pp19_w[42]), .i3(pp20_w[40]), .ci(stg1_co5[45]), .s(stg1_s5[46]), .c(stg1_c5[46]), .co(stg1_co5[46]));
counter_5to3 u_a15_47(.i0(pp17_w[47]), .i1(pp18_w[45]), .i2(pp19_w[43]), .i3(pp20_w[41]), .ci(stg1_co5[46]), .s(stg1_s5[47]), .c(stg1_c5[47]), .co(stg1_co5[47]));
counter_5to3 u_a15_48(.i0(pp17_w[48]), .i1(pp18_w[46]), .i2(pp19_w[44]), .i3(pp20_w[42]), .ci(stg1_co5[47]), .s(stg1_s5[48]), .c(stg1_c5[48]), .co(stg1_co5[48]));
counter_5to3 u_a15_49(.i0(pp17_w[49]), .i1(pp18_w[47]), .i2(pp19_w[45]), .i3(pp20_w[43]), .ci(stg1_co5[48]), .s(stg1_s5[49]), .c(stg1_c5[49]), .co(stg1_co5[49]));
counter_5to3 u_a15_50(.i0(pp17_w[50]), .i1(pp18_w[48]), .i2(pp19_w[46]), .i3(pp20_w[44]), .ci(stg1_co5[49]), .s(stg1_s5[50]), .c(stg1_c5[50]), .co(stg1_co5[50]));
counter_5to3 u_a15_51(.i0(pp17_w[51]), .i1(pp18_w[49]), .i2(pp19_w[47]), .i3(pp20_w[45]), .ci(stg1_co5[50]), .s(stg1_s5[51]), .c(stg1_c5[51]), .co(stg1_co5[51]));
counter_5to3 u_a15_52(.i0(pp17_w[52]), .i1(pp18_w[50]), .i2(pp19_w[48]), .i3(pp20_w[46]), .ci(stg1_co5[51]), .s(stg1_s5[52]), .c(stg1_c5[52]), .co(stg1_co5[52]));
counter_5to3 u_a15_53(.i0(pp17_w[53]), .i1(pp18_w[51]), .i2(pp19_w[49]), .i3(pp20_w[47]), .ci(stg1_co5[52]), .s(stg1_s5[53]), .c(stg1_c5[53]), .co(stg1_co5[53]));
counter_5to3 u_a15_54(.i0(pp17_w[54]), .i1(pp18_w[52]), .i2(pp19_w[50]), .i3(pp20_w[48]), .ci(stg1_co5[53]), .s(stg1_s5[54]), .c(stg1_c5[54]), .co(stg1_co5[54]));
counter_5to3 u_a15_55(.i0(pp17_w[55]), .i1(pp18_w[53]), .i2(pp19_w[51]), .i3(pp20_w[49]), .ci(stg1_co5[54]), .s(stg1_s5[55]), .c(stg1_c5[55]), .co(stg1_co5[55]));
counter_5to3 u_a15_56(.i0(pp17_w[56]), .i1(pp18_w[54]), .i2(pp19_w[52]), .i3(pp20_w[50]), .ci(stg1_co5[55]), .s(stg1_s5[56]), .c(stg1_c5[56]), .co(stg1_co5[56]));
counter_5to3 u_a15_57(.i0(pp17_w[57]), .i1(pp18_w[55]), .i2(pp19_w[53]), .i3(pp20_w[51]), .ci(stg1_co5[56]), .s(stg1_s5[57]), .c(stg1_c5[57]), .co(stg1_co5[57]));
counter_5to3 u_a15_58(.i0(pp17_w[58]), .i1(pp18_w[56]), .i2(pp19_w[54]), .i3(pp20_w[52]), .ci(stg1_co5[57]), .s(stg1_s5[58]), .c(stg1_c5[58]), .co(stg1_co5[58]));
counter_5to3 u_a15_59(.i0(pp17_w[59]), .i1(pp18_w[57]), .i2(pp19_w[55]), .i3(pp20_w[53]), .ci(stg1_co5[58]), .s(stg1_s5[59]), .c(stg1_c5[59]), .co(stg1_co5[59]));
counter_5to3 u_a15_60(.i0(pp17_w[60]), .i1(pp18_w[58]), .i2(pp19_w[56]), .i3(pp20_w[54]), .ci(stg1_co5[59]), .s(stg1_s5[60]), .c(stg1_c5[60]), .co(stg1_co5[60]));
counter_5to3 u_a15_61(.i0(pp17_w[61]), .i1(pp18_w[59]), .i2(pp19_w[57]), .i3(pp20_w[55]), .ci(stg1_co5[60]), .s(stg1_s5[61]), .c(stg1_c5[61]), .co(stg1_co5[61]));
counter_5to3 u_a15_62(.i0(pp17_w[62]), .i1(pp18_w[60]), .i2(pp19_w[58]), .i3(pp20_w[56]), .ci(stg1_co5[61]), .s(stg1_s5[62]), .c(stg1_c5[62]), .co(stg1_co5[62]));
counter_5to3 u_a15_63(.i0(pp17_w[63]), .i1(pp18_w[61]), .i2(pp19_w[59]), .i3(pp20_w[57]), .ci(stg1_co5[62]), .s(stg1_s5[63]), .c(stg1_c5[63]), .co(stg1_co5[63]));
counter_5to3 u_a15_64(.i0(pp17_w[64]), .i1(pp18_w[62]), .i2(pp19_w[60]), .i3(pp20_w[58]), .ci(stg1_co5[63]), .s(stg1_s5[64]), .c(stg1_c5[64]), .co(stg1_co5[64]));
counter_5to3 u_a15_65(.i0(pp17_w[65]), .i1(pp18_w[63]), .i2(pp19_w[61]), .i3(pp20_w[59]), .ci(stg1_co5[64]), .s(stg1_s5[65]), .c(stg1_c5[65]), .co(stg1_co5[65]));
counter_5to3 u_a15_66(.i0(pp17_w[65]), .i1(pp18_w[64]), .i2(pp19_w[62]), .i3(pp20_w[60]), .ci(stg1_co5[65]), .s(stg1_s5[66]), .c(stg1_c5[66]), .co(stg1_co5[66]));
counter_5to3 u_a15_67(.i0(pp17_w[65]), .i1(pp18_w[65]), .i2(pp19_w[63]), .i3(pp20_w[61]), .ci(stg1_co5[66]), .s(stg1_s5[67]), .c(stg1_c5[67]), .co(stg1_co5[67]));
counter_5to3 u_a15_68(.i0(pp17_w[65]), .i1(pp18_w[65]), .i2(pp19_w[64]), .i3(pp20_w[62]), .ci(stg1_co5[67]), .s(stg1_s5[68]), .c(stg1_c5[68]), .co(stg1_co5[68]));
counter_5to3 u_a15_69(.i0(pp17_w[65]), .i1(pp18_w[65]), .i2(pp19_w[65]), .i3(pp20_w[63]), .ci(stg1_co5[68]), .s(stg1_s5[69]), .c(stg1_c5[69]), .co(stg1_co5[69]));
counter_5to3 u_a15_70(.i0(pp17_w[65]), .i1(pp18_w[65]), .i2(pp19_w[65]), .i3(pp20_w[64]), .ci(stg1_co5[69]), .s(stg1_s5[70]), .c(stg1_c5[70]), .co(stg1_co5[70]));
counter_5to3 u_al5_71(.i0(pp17_w[65]), .i1(pp18_w[65]), .i2(pp19_w[65]), .i3(pp20_w[65]), .ci(stg1_co5[70]), .s(stg1_s5[71]), .c(stg1_c5[71]), .co(stg1_co5[71]));
counter_5to3 u_al5_72(.i0(pp17_w[65]), .i1(pp18_w[65]), .i2(pp19_w[65]), .i3(pp20_w[65]), .ci(stg1_co5[71]), .s(stg1_s5[72]), .c(stg1_c5[72]), .co(stg1_co5[72]));

// =========================== first stage 6th group ============================================================================================================
counter_5to3 u_a16_0 (.i0(pp21_w[0 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(1'b0        ), .s(stg1_s6[0 ]), .c(stg1_c6[0 ]), .co(stg1_co6[0 ]));
counter_5to3 u_a16_1 (.i0(pp21_w[1 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co6[0 ]), .s(stg1_s6[1 ]), .c(stg1_c6[1 ]), .co(stg1_co6[1 ]));
counter_5to3 u_a16_2 (.i0(pp21_w[2 ]), .i1(pp22_w[0 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co6[1 ]), .s(stg1_s6[2 ]), .c(stg1_c6[2 ]), .co(stg1_co6[2 ]));
counter_5to3 u_a16_3 (.i0(pp21_w[3 ]), .i1(pp22_w[1 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co6[2 ]), .s(stg1_s6[3 ]), .c(stg1_c6[3 ]), .co(stg1_co6[3 ]));
counter_5to3 u_a16_4 (.i0(pp21_w[4 ]), .i1(pp22_w[2 ]), .i2(pp23_w[0 ]), .i3(1'b0      ), .ci(stg1_co6[3 ]), .s(stg1_s6[4 ]), .c(stg1_c6[4 ]), .co(stg1_co6[4 ]));
counter_5to3 u_a16_5 (.i0(pp21_w[5 ]), .i1(pp22_w[3 ]), .i2(pp23_w[1 ]), .i3(1'b0      ), .ci(stg1_co6[4 ]), .s(stg1_s6[5 ]), .c(stg1_c6[5 ]), .co(stg1_co6[5 ]));
counter_5to3 u_a16_6 (.i0(pp21_w[6 ]), .i1(pp22_w[4 ]), .i2(pp23_w[2 ]), .i3(pp24_w[0 ]), .ci(stg1_co6[5 ]), .s(stg1_s6[6 ]), .c(stg1_c6[6 ]), .co(stg1_co6[6 ]));
counter_5to3 u_a16_7 (.i0(pp21_w[7 ]), .i1(pp22_w[5 ]), .i2(pp23_w[3 ]), .i3(pp24_w[1 ]), .ci(stg1_co6[6 ]), .s(stg1_s6[7 ]), .c(stg1_c6[7 ]), .co(stg1_co6[7 ]));
counter_5to3 u_a16_8 (.i0(pp21_w[8 ]), .i1(pp22_w[6 ]), .i2(pp23_w[4 ]), .i3(pp24_w[2 ]), .ci(stg1_co6[7 ]), .s(stg1_s6[8 ]), .c(stg1_c6[8 ]), .co(stg1_co6[8 ]));
counter_5to3 u_a16_9 (.i0(pp21_w[9 ]), .i1(pp22_w[7 ]), .i2(pp23_w[5 ]), .i3(pp24_w[3 ]), .ci(stg1_co6[8 ]), .s(stg1_s6[9 ]), .c(stg1_c6[9 ]), .co(stg1_co6[9 ]));
counter_5to3 u_a16_10(.i0(pp21_w[10]), .i1(pp22_w[8 ]), .i2(pp23_w[6 ]), .i3(pp24_w[4 ]), .ci(stg1_co6[9 ]), .s(stg1_s6[10]), .c(stg1_c6[10]), .co(stg1_co6[10]));
counter_5to3 u_a16_11(.i0(pp21_w[11]), .i1(pp22_w[9 ]), .i2(pp23_w[7 ]), .i3(pp24_w[5 ]), .ci(stg1_co6[10]), .s(stg1_s6[11]), .c(stg1_c6[11]), .co(stg1_co6[11]));
counter_5to3 u_a16_12(.i0(pp21_w[12]), .i1(pp22_w[10]), .i2(pp23_w[8 ]), .i3(pp24_w[6 ]), .ci(stg1_co6[11]), .s(stg1_s6[12]), .c(stg1_c6[12]), .co(stg1_co6[12]));
counter_5to3 u_a16_13(.i0(pp21_w[13]), .i1(pp22_w[11]), .i2(pp23_w[9 ]), .i3(pp24_w[7 ]), .ci(stg1_co6[12]), .s(stg1_s6[13]), .c(stg1_c6[13]), .co(stg1_co6[13]));
counter_5to3 u_a16_14(.i0(pp21_w[14]), .i1(pp22_w[12]), .i2(pp23_w[10]), .i3(pp24_w[8 ]), .ci(stg1_co6[13]), .s(stg1_s6[14]), .c(stg1_c6[14]), .co(stg1_co6[14]));
counter_5to3 u_a16_15(.i0(pp21_w[15]), .i1(pp22_w[13]), .i2(pp23_w[11]), .i3(pp24_w[9 ]), .ci(stg1_co6[14]), .s(stg1_s6[15]), .c(stg1_c6[15]), .co(stg1_co6[15]));
counter_5to3 u_a16_16(.i0(pp21_w[16]), .i1(pp22_w[14]), .i2(pp23_w[12]), .i3(pp24_w[10]), .ci(stg1_co6[15]), .s(stg1_s6[16]), .c(stg1_c6[16]), .co(stg1_co6[16]));
counter_5to3 u_a16_17(.i0(pp21_w[17]), .i1(pp22_w[15]), .i2(pp23_w[13]), .i3(pp24_w[11]), .ci(stg1_co6[16]), .s(stg1_s6[17]), .c(stg1_c6[17]), .co(stg1_co6[17]));
counter_5to3 u_a16_18(.i0(pp21_w[18]), .i1(pp22_w[16]), .i2(pp23_w[14]), .i3(pp24_w[12]), .ci(stg1_co6[17]), .s(stg1_s6[18]), .c(stg1_c6[18]), .co(stg1_co6[18]));
counter_5to3 u_a16_19(.i0(pp21_w[19]), .i1(pp22_w[17]), .i2(pp23_w[15]), .i3(pp24_w[13]), .ci(stg1_co6[18]), .s(stg1_s6[19]), .c(stg1_c6[19]), .co(stg1_co6[19]));
counter_5to3 u_a16_20(.i0(pp21_w[20]), .i1(pp22_w[18]), .i2(pp23_w[16]), .i3(pp24_w[14]), .ci(stg1_co6[19]), .s(stg1_s6[20]), .c(stg1_c6[20]), .co(stg1_co6[20]));
counter_5to3 u_a16_21(.i0(pp21_w[21]), .i1(pp22_w[19]), .i2(pp23_w[17]), .i3(pp24_w[15]), .ci(stg1_co6[20]), .s(stg1_s6[21]), .c(stg1_c6[21]), .co(stg1_co6[21]));
counter_5to3 u_a16_22(.i0(pp21_w[22]), .i1(pp22_w[20]), .i2(pp23_w[18]), .i3(pp24_w[16]), .ci(stg1_co6[21]), .s(stg1_s6[22]), .c(stg1_c6[22]), .co(stg1_co6[22]));
counter_5to3 u_a16_23(.i0(pp21_w[23]), .i1(pp22_w[21]), .i2(pp23_w[19]), .i3(pp24_w[17]), .ci(stg1_co6[22]), .s(stg1_s6[23]), .c(stg1_c6[23]), .co(stg1_co6[23]));
counter_5to3 u_a16_24(.i0(pp21_w[24]), .i1(pp22_w[22]), .i2(pp23_w[20]), .i3(pp24_w[18]), .ci(stg1_co6[23]), .s(stg1_s6[24]), .c(stg1_c6[24]), .co(stg1_co6[24]));
counter_5to3 u_a16_25(.i0(pp21_w[25]), .i1(pp22_w[23]), .i2(pp23_w[21]), .i3(pp24_w[19]), .ci(stg1_co6[24]), .s(stg1_s6[25]), .c(stg1_c6[25]), .co(stg1_co6[25]));
counter_5to3 u_a16_26(.i0(pp21_w[26]), .i1(pp22_w[24]), .i2(pp23_w[22]), .i3(pp24_w[20]), .ci(stg1_co6[25]), .s(stg1_s6[26]), .c(stg1_c6[26]), .co(stg1_co6[26]));
counter_5to3 u_a16_27(.i0(pp21_w[27]), .i1(pp22_w[25]), .i2(pp23_w[23]), .i3(pp24_w[21]), .ci(stg1_co6[26]), .s(stg1_s6[27]), .c(stg1_c6[27]), .co(stg1_co6[27]));
counter_5to3 u_a16_28(.i0(pp21_w[28]), .i1(pp22_w[26]), .i2(pp23_w[24]), .i3(pp24_w[22]), .ci(stg1_co6[27]), .s(stg1_s6[28]), .c(stg1_c6[28]), .co(stg1_co6[28]));
counter_5to3 u_a16_29(.i0(pp21_w[29]), .i1(pp22_w[27]), .i2(pp23_w[25]), .i3(pp24_w[23]), .ci(stg1_co6[28]), .s(stg1_s6[29]), .c(stg1_c6[29]), .co(stg1_co6[29]));
counter_5to3 u_a16_30(.i0(pp21_w[30]), .i1(pp22_w[28]), .i2(pp23_w[26]), .i3(pp24_w[24]), .ci(stg1_co6[29]), .s(stg1_s6[30]), .c(stg1_c6[30]), .co(stg1_co6[30]));
counter_5to3 u_a16_31(.i0(pp21_w[31]), .i1(pp22_w[29]), .i2(pp23_w[27]), .i3(pp24_w[25]), .ci(stg1_co6[30]), .s(stg1_s6[31]), .c(stg1_c6[31]), .co(stg1_co6[31]));
counter_5to3 u_a16_32(.i0(pp21_w[32]), .i1(pp22_w[30]), .i2(pp23_w[28]), .i3(pp24_w[26]), .ci(stg1_co6[31]), .s(stg1_s6[32]), .c(stg1_c6[32]), .co(stg1_co6[32]));
counter_5to3 u_a16_33(.i0(pp21_w[33]), .i1(pp22_w[31]), .i2(pp23_w[29]), .i3(pp24_w[27]), .ci(stg1_co6[32]), .s(stg1_s6[33]), .c(stg1_c6[33]), .co(stg1_co6[33]));
counter_5to3 u_a16_34(.i0(pp21_w[34]), .i1(pp22_w[32]), .i2(pp23_w[30]), .i3(pp24_w[28]), .ci(stg1_co6[33]), .s(stg1_s6[34]), .c(stg1_c6[34]), .co(stg1_co6[34]));
counter_5to3 u_a16_35(.i0(pp21_w[35]), .i1(pp22_w[33]), .i2(pp23_w[31]), .i3(pp24_w[29]), .ci(stg1_co6[34]), .s(stg1_s6[35]), .c(stg1_c6[35]), .co(stg1_co6[35]));
counter_5to3 u_a16_36(.i0(pp21_w[36]), .i1(pp22_w[34]), .i2(pp23_w[32]), .i3(pp24_w[30]), .ci(stg1_co6[35]), .s(stg1_s6[36]), .c(stg1_c6[36]), .co(stg1_co6[36]));
counter_5to3 u_a16_37(.i0(pp21_w[37]), .i1(pp22_w[35]), .i2(pp23_w[33]), .i3(pp24_w[31]), .ci(stg1_co6[36]), .s(stg1_s6[37]), .c(stg1_c6[37]), .co(stg1_co6[37]));
counter_5to3 u_a16_38(.i0(pp21_w[38]), .i1(pp22_w[36]), .i2(pp23_w[34]), .i3(pp24_w[32]), .ci(stg1_co6[37]), .s(stg1_s6[38]), .c(stg1_c6[38]), .co(stg1_co6[38]));
counter_5to3 u_a16_39(.i0(pp21_w[39]), .i1(pp22_w[37]), .i2(pp23_w[35]), .i3(pp24_w[33]), .ci(stg1_co6[38]), .s(stg1_s6[39]), .c(stg1_c6[39]), .co(stg1_co6[39]));
counter_5to3 u_a16_40(.i0(pp21_w[40]), .i1(pp22_w[38]), .i2(pp23_w[36]), .i3(pp24_w[34]), .ci(stg1_co6[39]), .s(stg1_s6[40]), .c(stg1_c6[40]), .co(stg1_co6[40]));
counter_5to3 u_a16_41(.i0(pp21_w[41]), .i1(pp22_w[39]), .i2(pp23_w[37]), .i3(pp24_w[35]), .ci(stg1_co6[40]), .s(stg1_s6[41]), .c(stg1_c6[41]), .co(stg1_co6[41]));
counter_5to3 u_a16_42(.i0(pp21_w[42]), .i1(pp22_w[40]), .i2(pp23_w[38]), .i3(pp24_w[36]), .ci(stg1_co6[41]), .s(stg1_s6[42]), .c(stg1_c6[42]), .co(stg1_co6[42]));
counter_5to3 u_a16_43(.i0(pp21_w[43]), .i1(pp22_w[41]), .i2(pp23_w[39]), .i3(pp24_w[37]), .ci(stg1_co6[42]), .s(stg1_s6[43]), .c(stg1_c6[43]), .co(stg1_co6[43]));
counter_5to3 u_a16_44(.i0(pp21_w[44]), .i1(pp22_w[42]), .i2(pp23_w[40]), .i3(pp24_w[38]), .ci(stg1_co6[43]), .s(stg1_s6[44]), .c(stg1_c6[44]), .co(stg1_co6[44]));
counter_5to3 u_a16_45(.i0(pp21_w[45]), .i1(pp22_w[43]), .i2(pp23_w[41]), .i3(pp24_w[39]), .ci(stg1_co6[44]), .s(stg1_s6[45]), .c(stg1_c6[45]), .co(stg1_co6[45]));
counter_5to3 u_a16_46(.i0(pp21_w[46]), .i1(pp22_w[44]), .i2(pp23_w[42]), .i3(pp24_w[40]), .ci(stg1_co6[45]), .s(stg1_s6[46]), .c(stg1_c6[46]), .co(stg1_co6[46]));
counter_5to3 u_a16_47(.i0(pp21_w[47]), .i1(pp22_w[45]), .i2(pp23_w[43]), .i3(pp24_w[41]), .ci(stg1_co6[46]), .s(stg1_s6[47]), .c(stg1_c6[47]), .co(stg1_co6[47]));
counter_5to3 u_a16_48(.i0(pp21_w[48]), .i1(pp22_w[46]), .i2(pp23_w[44]), .i3(pp24_w[42]), .ci(stg1_co6[47]), .s(stg1_s6[48]), .c(stg1_c6[48]), .co(stg1_co6[48]));
counter_5to3 u_a16_49(.i0(pp21_w[49]), .i1(pp22_w[47]), .i2(pp23_w[45]), .i3(pp24_w[43]), .ci(stg1_co6[48]), .s(stg1_s6[49]), .c(stg1_c6[49]), .co(stg1_co6[49]));
counter_5to3 u_a16_50(.i0(pp21_w[50]), .i1(pp22_w[48]), .i2(pp23_w[46]), .i3(pp24_w[44]), .ci(stg1_co6[49]), .s(stg1_s6[50]), .c(stg1_c6[50]), .co(stg1_co6[50]));
counter_5to3 u_a16_51(.i0(pp21_w[51]), .i1(pp22_w[49]), .i2(pp23_w[47]), .i3(pp24_w[45]), .ci(stg1_co6[50]), .s(stg1_s6[51]), .c(stg1_c6[51]), .co(stg1_co6[51]));
counter_5to3 u_a16_52(.i0(pp21_w[52]), .i1(pp22_w[50]), .i2(pp23_w[48]), .i3(pp24_w[46]), .ci(stg1_co6[51]), .s(stg1_s6[52]), .c(stg1_c6[52]), .co(stg1_co6[52]));
counter_5to3 u_a16_53(.i0(pp21_w[53]), .i1(pp22_w[51]), .i2(pp23_w[49]), .i3(pp24_w[47]), .ci(stg1_co6[52]), .s(stg1_s6[53]), .c(stg1_c6[53]), .co(stg1_co6[53]));
counter_5to3 u_a16_54(.i0(pp21_w[54]), .i1(pp22_w[52]), .i2(pp23_w[50]), .i3(pp24_w[48]), .ci(stg1_co6[53]), .s(stg1_s6[54]), .c(stg1_c6[54]), .co(stg1_co6[54]));
counter_5to3 u_a16_55(.i0(pp21_w[55]), .i1(pp22_w[53]), .i2(pp23_w[51]), .i3(pp24_w[49]), .ci(stg1_co6[54]), .s(stg1_s6[55]), .c(stg1_c6[55]), .co(stg1_co6[55]));
counter_5to3 u_a16_56(.i0(pp21_w[56]), .i1(pp22_w[54]), .i2(pp23_w[52]), .i3(pp24_w[50]), .ci(stg1_co6[55]), .s(stg1_s6[56]), .c(stg1_c6[56]), .co(stg1_co6[56]));
counter_5to3 u_a16_57(.i0(pp21_w[57]), .i1(pp22_w[55]), .i2(pp23_w[53]), .i3(pp24_w[51]), .ci(stg1_co6[56]), .s(stg1_s6[57]), .c(stg1_c6[57]), .co(stg1_co6[57]));
counter_5to3 u_a16_58(.i0(pp21_w[58]), .i1(pp22_w[56]), .i2(pp23_w[54]), .i3(pp24_w[52]), .ci(stg1_co6[57]), .s(stg1_s6[58]), .c(stg1_c6[58]), .co(stg1_co6[58]));
counter_5to3 u_a16_59(.i0(pp21_w[59]), .i1(pp22_w[57]), .i2(pp23_w[55]), .i3(pp24_w[53]), .ci(stg1_co6[58]), .s(stg1_s6[59]), .c(stg1_c6[59]), .co(stg1_co6[59]));
counter_5to3 u_a16_60(.i0(pp21_w[60]), .i1(pp22_w[58]), .i2(pp23_w[56]), .i3(pp24_w[54]), .ci(stg1_co6[59]), .s(stg1_s6[60]), .c(stg1_c6[60]), .co(stg1_co6[60]));
counter_5to3 u_a16_61(.i0(pp21_w[61]), .i1(pp22_w[59]), .i2(pp23_w[57]), .i3(pp24_w[55]), .ci(stg1_co6[60]), .s(stg1_s6[61]), .c(stg1_c6[61]), .co(stg1_co6[61]));
counter_5to3 u_a16_62(.i0(pp21_w[62]), .i1(pp22_w[60]), .i2(pp23_w[58]), .i3(pp24_w[56]), .ci(stg1_co6[61]), .s(stg1_s6[62]), .c(stg1_c6[62]), .co(stg1_co6[62]));
counter_5to3 u_a16_63(.i0(pp21_w[63]), .i1(pp22_w[61]), .i2(pp23_w[59]), .i3(pp24_w[57]), .ci(stg1_co6[62]), .s(stg1_s6[63]), .c(stg1_c6[63]), .co(stg1_co6[63]));
counter_5to3 u_a16_64(.i0(pp21_w[64]), .i1(pp22_w[62]), .i2(pp23_w[60]), .i3(pp24_w[58]), .ci(stg1_co6[63]), .s(stg1_s6[64]), .c(stg1_c6[64]), .co(stg1_co6[64]));
counter_5to3 u_a16_65(.i0(pp21_w[65]), .i1(pp22_w[63]), .i2(pp23_w[61]), .i3(pp24_w[59]), .ci(stg1_co6[64]), .s(stg1_s6[65]), .c(stg1_c6[65]), .co(stg1_co6[65]));
counter_5to3 u_a16_66(.i0(pp21_w[65]), .i1(pp22_w[64]), .i2(pp23_w[62]), .i3(pp24_w[60]), .ci(stg1_co6[65]), .s(stg1_s6[66]), .c(stg1_c6[66]), .co(stg1_co6[66]));
counter_5to3 u_a16_67(.i0(pp21_w[65]), .i1(pp22_w[65]), .i2(pp23_w[63]), .i3(pp24_w[61]), .ci(stg1_co6[66]), .s(stg1_s6[67]), .c(stg1_c6[67]), .co(stg1_co6[67]));
counter_5to3 u_a16_68(.i0(pp21_w[65]), .i1(pp22_w[65]), .i2(pp23_w[64]), .i3(pp24_w[62]), .ci(stg1_co6[67]), .s(stg1_s6[68]), .c(stg1_c6[68]), .co(stg1_co6[68]));
counter_5to3 u_a16_69(.i0(pp21_w[65]), .i1(pp22_w[65]), .i2(pp23_w[65]), .i3(pp24_w[63]), .ci(stg1_co6[68]), .s(stg1_s6[69]), .c(stg1_c6[69]), .co(stg1_co6[69]));
counter_5to3 u_a16_70(.i0(pp21_w[65]), .i1(pp22_w[65]), .i2(pp23_w[65]), .i3(pp24_w[64]), .ci(stg1_co6[69]), .s(stg1_s6[70]), .c(stg1_c6[70]), .co(stg1_co6[70]));
counter_5to3 u_al6_71(.i0(pp21_w[65]), .i1(pp22_w[65]), .i2(pp23_w[65]), .i3(pp24_w[65]), .ci(stg1_co6[70]), .s(stg1_s6[71]), .c(stg1_c6[71]), .co(stg1_co6[71]));
counter_5to3 u_al6_72(.i0(pp21_w[65]), .i1(pp22_w[65]), .i2(pp23_w[65]), .i3(pp24_w[65]), .ci(stg1_co6[71]), .s(stg1_s6[72]), .c(stg1_c6[72]), .co(stg1_co6[72]));

// =========================== first stage 7th group ============================================================================================================
counter_5to3 u_a17_0 (.i0(pp25_w[0 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(1'b0        ), .s(stg1_s7[0 ]), .c(stg1_c7[0 ]), .co(stg1_co7[0 ]));
counter_5to3 u_a17_1 (.i0(pp25_w[1 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co7[0 ]), .s(stg1_s7[1 ]), .c(stg1_c7[1 ]), .co(stg1_co7[1 ]));
counter_5to3 u_a17_2 (.i0(pp25_w[2 ]), .i1(pp26_w[0 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co7[1 ]), .s(stg1_s7[2 ]), .c(stg1_c7[2 ]), .co(stg1_co7[2 ]));
counter_5to3 u_a17_3 (.i0(pp25_w[3 ]), .i1(pp26_w[1 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co7[2 ]), .s(stg1_s7[3 ]), .c(stg1_c7[3 ]), .co(stg1_co7[3 ]));
counter_5to3 u_a17_4 (.i0(pp25_w[4 ]), .i1(pp26_w[2 ]), .i2(pp27_w[0 ]), .i3(1'b0      ), .ci(stg1_co7[3 ]), .s(stg1_s7[4 ]), .c(stg1_c7[4 ]), .co(stg1_co7[4 ]));
counter_5to3 u_a17_5 (.i0(pp25_w[5 ]), .i1(pp26_w[3 ]), .i2(pp27_w[1 ]), .i3(1'b0      ), .ci(stg1_co7[4 ]), .s(stg1_s7[5 ]), .c(stg1_c7[5 ]), .co(stg1_co7[5 ]));
counter_5to3 u_a17_6 (.i0(pp25_w[6 ]), .i1(pp26_w[4 ]), .i2(pp27_w[2 ]), .i3(pp28_w[0 ]), .ci(stg1_co7[5 ]), .s(stg1_s7[6 ]), .c(stg1_c7[6 ]), .co(stg1_co7[6 ]));
counter_5to3 u_a17_7 (.i0(pp25_w[7 ]), .i1(pp26_w[5 ]), .i2(pp27_w[3 ]), .i3(pp28_w[1 ]), .ci(stg1_co7[6 ]), .s(stg1_s7[7 ]), .c(stg1_c7[7 ]), .co(stg1_co7[7 ]));
counter_5to3 u_a17_8 (.i0(pp25_w[8 ]), .i1(pp26_w[6 ]), .i2(pp27_w[4 ]), .i3(pp28_w[2 ]), .ci(stg1_co7[7 ]), .s(stg1_s7[8 ]), .c(stg1_c7[8 ]), .co(stg1_co7[8 ]));
counter_5to3 u_a17_9 (.i0(pp25_w[9 ]), .i1(pp26_w[7 ]), .i2(pp27_w[5 ]), .i3(pp28_w[3 ]), .ci(stg1_co7[8 ]), .s(stg1_s7[9 ]), .c(stg1_c7[9 ]), .co(stg1_co7[9 ]));
counter_5to3 u_a17_10(.i0(pp25_w[10]), .i1(pp26_w[8 ]), .i2(pp27_w[6 ]), .i3(pp28_w[4 ]), .ci(stg1_co7[9 ]), .s(stg1_s7[10]), .c(stg1_c7[10]), .co(stg1_co7[10]));
counter_5to3 u_a17_11(.i0(pp25_w[11]), .i1(pp26_w[9 ]), .i2(pp27_w[7 ]), .i3(pp28_w[5 ]), .ci(stg1_co7[10]), .s(stg1_s7[11]), .c(stg1_c7[11]), .co(stg1_co7[11]));
counter_5to3 u_a17_12(.i0(pp25_w[12]), .i1(pp26_w[10]), .i2(pp27_w[8 ]), .i3(pp28_w[6 ]), .ci(stg1_co7[11]), .s(stg1_s7[12]), .c(stg1_c7[12]), .co(stg1_co7[12]));
counter_5to3 u_a17_13(.i0(pp25_w[13]), .i1(pp26_w[11]), .i2(pp27_w[9 ]), .i3(pp28_w[7 ]), .ci(stg1_co7[12]), .s(stg1_s7[13]), .c(stg1_c7[13]), .co(stg1_co7[13]));
counter_5to3 u_a17_14(.i0(pp25_w[14]), .i1(pp26_w[12]), .i2(pp27_w[10]), .i3(pp28_w[8 ]), .ci(stg1_co7[13]), .s(stg1_s7[14]), .c(stg1_c7[14]), .co(stg1_co7[14]));
counter_5to3 u_a17_15(.i0(pp25_w[15]), .i1(pp26_w[13]), .i2(pp27_w[11]), .i3(pp28_w[9 ]), .ci(stg1_co7[14]), .s(stg1_s7[15]), .c(stg1_c7[15]), .co(stg1_co7[15]));
counter_5to3 u_a17_16(.i0(pp25_w[16]), .i1(pp26_w[14]), .i2(pp27_w[12]), .i3(pp28_w[10]), .ci(stg1_co7[15]), .s(stg1_s7[16]), .c(stg1_c7[16]), .co(stg1_co7[16]));
counter_5to3 u_a17_17(.i0(pp25_w[17]), .i1(pp26_w[15]), .i2(pp27_w[13]), .i3(pp28_w[11]), .ci(stg1_co7[16]), .s(stg1_s7[17]), .c(stg1_c7[17]), .co(stg1_co7[17]));
counter_5to3 u_a17_18(.i0(pp25_w[18]), .i1(pp26_w[16]), .i2(pp27_w[14]), .i3(pp28_w[12]), .ci(stg1_co7[17]), .s(stg1_s7[18]), .c(stg1_c7[18]), .co(stg1_co7[18]));
counter_5to3 u_a17_19(.i0(pp25_w[19]), .i1(pp26_w[17]), .i2(pp27_w[15]), .i3(pp28_w[13]), .ci(stg1_co7[18]), .s(stg1_s7[19]), .c(stg1_c7[19]), .co(stg1_co7[19]));
counter_5to3 u_a17_20(.i0(pp25_w[20]), .i1(pp26_w[18]), .i2(pp27_w[16]), .i3(pp28_w[14]), .ci(stg1_co7[19]), .s(stg1_s7[20]), .c(stg1_c7[20]), .co(stg1_co7[20]));
counter_5to3 u_a17_21(.i0(pp25_w[21]), .i1(pp26_w[19]), .i2(pp27_w[17]), .i3(pp28_w[15]), .ci(stg1_co7[20]), .s(stg1_s7[21]), .c(stg1_c7[21]), .co(stg1_co7[21]));
counter_5to3 u_a17_22(.i0(pp25_w[22]), .i1(pp26_w[20]), .i2(pp27_w[18]), .i3(pp28_w[16]), .ci(stg1_co7[21]), .s(stg1_s7[22]), .c(stg1_c7[22]), .co(stg1_co7[22]));
counter_5to3 u_a17_23(.i0(pp25_w[23]), .i1(pp26_w[21]), .i2(pp27_w[19]), .i3(pp28_w[17]), .ci(stg1_co7[22]), .s(stg1_s7[23]), .c(stg1_c7[23]), .co(stg1_co7[23]));
counter_5to3 u_a17_24(.i0(pp25_w[24]), .i1(pp26_w[22]), .i2(pp27_w[20]), .i3(pp28_w[18]), .ci(stg1_co7[23]), .s(stg1_s7[24]), .c(stg1_c7[24]), .co(stg1_co7[24]));
counter_5to3 u_a17_25(.i0(pp25_w[25]), .i1(pp26_w[23]), .i2(pp27_w[21]), .i3(pp28_w[19]), .ci(stg1_co7[24]), .s(stg1_s7[25]), .c(stg1_c7[25]), .co(stg1_co7[25]));
counter_5to3 u_a17_26(.i0(pp25_w[26]), .i1(pp26_w[24]), .i2(pp27_w[22]), .i3(pp28_w[20]), .ci(stg1_co7[25]), .s(stg1_s7[26]), .c(stg1_c7[26]), .co(stg1_co7[26]));
counter_5to3 u_a17_27(.i0(pp25_w[27]), .i1(pp26_w[25]), .i2(pp27_w[23]), .i3(pp28_w[21]), .ci(stg1_co7[26]), .s(stg1_s7[27]), .c(stg1_c7[27]), .co(stg1_co7[27]));
counter_5to3 u_a17_28(.i0(pp25_w[28]), .i1(pp26_w[26]), .i2(pp27_w[24]), .i3(pp28_w[22]), .ci(stg1_co7[27]), .s(stg1_s7[28]), .c(stg1_c7[28]), .co(stg1_co7[28]));
counter_5to3 u_a17_29(.i0(pp25_w[29]), .i1(pp26_w[27]), .i2(pp27_w[25]), .i3(pp28_w[23]), .ci(stg1_co7[28]), .s(stg1_s7[29]), .c(stg1_c7[29]), .co(stg1_co7[29]));
counter_5to3 u_a17_30(.i0(pp25_w[30]), .i1(pp26_w[28]), .i2(pp27_w[26]), .i3(pp28_w[24]), .ci(stg1_co7[29]), .s(stg1_s7[30]), .c(stg1_c7[30]), .co(stg1_co7[30]));
counter_5to3 u_a17_31(.i0(pp25_w[31]), .i1(pp26_w[29]), .i2(pp27_w[27]), .i3(pp28_w[25]), .ci(stg1_co7[30]), .s(stg1_s7[31]), .c(stg1_c7[31]), .co(stg1_co7[31]));
counter_5to3 u_a17_32(.i0(pp25_w[32]), .i1(pp26_w[30]), .i2(pp27_w[28]), .i3(pp28_w[26]), .ci(stg1_co7[31]), .s(stg1_s7[32]), .c(stg1_c7[32]), .co(stg1_co7[32]));
counter_5to3 u_a17_33(.i0(pp25_w[33]), .i1(pp26_w[31]), .i2(pp27_w[29]), .i3(pp28_w[27]), .ci(stg1_co7[32]), .s(stg1_s7[33]), .c(stg1_c7[33]), .co(stg1_co7[33]));
counter_5to3 u_a17_34(.i0(pp25_w[34]), .i1(pp26_w[32]), .i2(pp27_w[30]), .i3(pp28_w[28]), .ci(stg1_co7[33]), .s(stg1_s7[34]), .c(stg1_c7[34]), .co(stg1_co7[34]));
counter_5to3 u_a17_35(.i0(pp25_w[35]), .i1(pp26_w[33]), .i2(pp27_w[31]), .i3(pp28_w[29]), .ci(stg1_co7[34]), .s(stg1_s7[35]), .c(stg1_c7[35]), .co(stg1_co7[35]));
counter_5to3 u_a17_36(.i0(pp25_w[36]), .i1(pp26_w[34]), .i2(pp27_w[32]), .i3(pp28_w[30]), .ci(stg1_co7[35]), .s(stg1_s7[36]), .c(stg1_c7[36]), .co(stg1_co7[36]));
counter_5to3 u_a17_37(.i0(pp25_w[37]), .i1(pp26_w[35]), .i2(pp27_w[33]), .i3(pp28_w[31]), .ci(stg1_co7[36]), .s(stg1_s7[37]), .c(stg1_c7[37]), .co(stg1_co7[37]));
counter_5to3 u_a17_38(.i0(pp25_w[38]), .i1(pp26_w[36]), .i2(pp27_w[34]), .i3(pp28_w[32]), .ci(stg1_co7[37]), .s(stg1_s7[38]), .c(stg1_c7[38]), .co(stg1_co7[38]));
counter_5to3 u_a17_39(.i0(pp25_w[39]), .i1(pp26_w[37]), .i2(pp27_w[35]), .i3(pp28_w[33]), .ci(stg1_co7[38]), .s(stg1_s7[39]), .c(stg1_c7[39]), .co(stg1_co7[39]));
counter_5to3 u_a17_40(.i0(pp25_w[40]), .i1(pp26_w[38]), .i2(pp27_w[36]), .i3(pp28_w[34]), .ci(stg1_co7[39]), .s(stg1_s7[40]), .c(stg1_c7[40]), .co(stg1_co7[40]));
counter_5to3 u_a17_41(.i0(pp25_w[41]), .i1(pp26_w[39]), .i2(pp27_w[37]), .i3(pp28_w[35]), .ci(stg1_co7[40]), .s(stg1_s7[41]), .c(stg1_c7[41]), .co(stg1_co7[41]));
counter_5to3 u_a17_42(.i0(pp25_w[42]), .i1(pp26_w[40]), .i2(pp27_w[38]), .i3(pp28_w[36]), .ci(stg1_co7[41]), .s(stg1_s7[42]), .c(stg1_c7[42]), .co(stg1_co7[42]));
counter_5to3 u_a17_43(.i0(pp25_w[43]), .i1(pp26_w[41]), .i2(pp27_w[39]), .i3(pp28_w[37]), .ci(stg1_co7[42]), .s(stg1_s7[43]), .c(stg1_c7[43]), .co(stg1_co7[43]));
counter_5to3 u_a17_44(.i0(pp25_w[44]), .i1(pp26_w[42]), .i2(pp27_w[40]), .i3(pp28_w[38]), .ci(stg1_co7[43]), .s(stg1_s7[44]), .c(stg1_c7[44]), .co(stg1_co7[44]));
counter_5to3 u_a17_45(.i0(pp25_w[45]), .i1(pp26_w[43]), .i2(pp27_w[41]), .i3(pp28_w[39]), .ci(stg1_co7[44]), .s(stg1_s7[45]), .c(stg1_c7[45]), .co(stg1_co7[45]));
counter_5to3 u_a17_46(.i0(pp25_w[46]), .i1(pp26_w[44]), .i2(pp27_w[42]), .i3(pp28_w[40]), .ci(stg1_co7[45]), .s(stg1_s7[46]), .c(stg1_c7[46]), .co(stg1_co7[46]));
counter_5to3 u_a17_47(.i0(pp25_w[47]), .i1(pp26_w[45]), .i2(pp27_w[43]), .i3(pp28_w[41]), .ci(stg1_co7[46]), .s(stg1_s7[47]), .c(stg1_c7[47]), .co(stg1_co7[47]));
counter_5to3 u_a17_48(.i0(pp25_w[48]), .i1(pp26_w[46]), .i2(pp27_w[44]), .i3(pp28_w[42]), .ci(stg1_co7[47]), .s(stg1_s7[48]), .c(stg1_c7[48]), .co(stg1_co7[48]));
counter_5to3 u_a17_49(.i0(pp25_w[49]), .i1(pp26_w[47]), .i2(pp27_w[45]), .i3(pp28_w[43]), .ci(stg1_co7[48]), .s(stg1_s7[49]), .c(stg1_c7[49]), .co(stg1_co7[49]));
counter_5to3 u_a17_50(.i0(pp25_w[50]), .i1(pp26_w[48]), .i2(pp27_w[46]), .i3(pp28_w[44]), .ci(stg1_co7[49]), .s(stg1_s7[50]), .c(stg1_c7[50]), .co(stg1_co7[50]));
counter_5to3 u_a17_51(.i0(pp25_w[51]), .i1(pp26_w[49]), .i2(pp27_w[47]), .i3(pp28_w[45]), .ci(stg1_co7[50]), .s(stg1_s7[51]), .c(stg1_c7[51]), .co(stg1_co7[51]));
counter_5to3 u_a17_52(.i0(pp25_w[52]), .i1(pp26_w[50]), .i2(pp27_w[48]), .i3(pp28_w[46]), .ci(stg1_co7[51]), .s(stg1_s7[52]), .c(stg1_c7[52]), .co(stg1_co7[52]));
counter_5to3 u_a17_53(.i0(pp25_w[53]), .i1(pp26_w[51]), .i2(pp27_w[49]), .i3(pp28_w[47]), .ci(stg1_co7[52]), .s(stg1_s7[53]), .c(stg1_c7[53]), .co(stg1_co7[53]));
counter_5to3 u_a17_54(.i0(pp25_w[54]), .i1(pp26_w[52]), .i2(pp27_w[50]), .i3(pp28_w[48]), .ci(stg1_co7[53]), .s(stg1_s7[54]), .c(stg1_c7[54]), .co(stg1_co7[54]));
counter_5to3 u_a17_55(.i0(pp25_w[55]), .i1(pp26_w[53]), .i2(pp27_w[51]), .i3(pp28_w[49]), .ci(stg1_co7[54]), .s(stg1_s7[55]), .c(stg1_c7[55]), .co(stg1_co7[55]));
counter_5to3 u_a17_56(.i0(pp25_w[56]), .i1(pp26_w[54]), .i2(pp27_w[52]), .i3(pp28_w[50]), .ci(stg1_co7[55]), .s(stg1_s7[56]), .c(stg1_c7[56]), .co(stg1_co7[56]));
counter_5to3 u_a17_57(.i0(pp25_w[57]), .i1(pp26_w[55]), .i2(pp27_w[53]), .i3(pp28_w[51]), .ci(stg1_co7[56]), .s(stg1_s7[57]), .c(stg1_c7[57]), .co(stg1_co7[57]));
counter_5to3 u_a17_58(.i0(pp25_w[58]), .i1(pp26_w[56]), .i2(pp27_w[54]), .i3(pp28_w[52]), .ci(stg1_co7[57]), .s(stg1_s7[58]), .c(stg1_c7[58]), .co(stg1_co7[58]));
counter_5to3 u_a17_59(.i0(pp25_w[59]), .i1(pp26_w[57]), .i2(pp27_w[55]), .i3(pp28_w[53]), .ci(stg1_co7[58]), .s(stg1_s7[59]), .c(stg1_c7[59]), .co(stg1_co7[59]));
counter_5to3 u_a17_60(.i0(pp25_w[60]), .i1(pp26_w[58]), .i2(pp27_w[56]), .i3(pp28_w[54]), .ci(stg1_co7[59]), .s(stg1_s7[60]), .c(stg1_c7[60]), .co(stg1_co7[60]));
counter_5to3 u_a17_61(.i0(pp25_w[61]), .i1(pp26_w[59]), .i2(pp27_w[57]), .i3(pp28_w[55]), .ci(stg1_co7[60]), .s(stg1_s7[61]), .c(stg1_c7[61]), .co(stg1_co7[61]));
counter_5to3 u_a17_62(.i0(pp25_w[62]), .i1(pp26_w[60]), .i2(pp27_w[58]), .i3(pp28_w[56]), .ci(stg1_co7[61]), .s(stg1_s7[62]), .c(stg1_c7[62]), .co(stg1_co7[62]));
counter_5to3 u_a17_63(.i0(pp25_w[63]), .i1(pp26_w[61]), .i2(pp27_w[59]), .i3(pp28_w[57]), .ci(stg1_co7[62]), .s(stg1_s7[63]), .c(stg1_c7[63]), .co(stg1_co7[63]));
counter_5to3 u_a17_64(.i0(pp25_w[64]), .i1(pp26_w[62]), .i2(pp27_w[60]), .i3(pp28_w[58]), .ci(stg1_co7[63]), .s(stg1_s7[64]), .c(stg1_c7[64]), .co(stg1_co7[64]));
counter_5to3 u_a17_65(.i0(pp25_w[65]), .i1(pp26_w[63]), .i2(pp27_w[61]), .i3(pp28_w[59]), .ci(stg1_co7[64]), .s(stg1_s7[65]), .c(stg1_c7[65]), .co(stg1_co7[65]));
counter_5to3 u_a17_66(.i0(pp25_w[65]), .i1(pp26_w[64]), .i2(pp27_w[62]), .i3(pp28_w[60]), .ci(stg1_co7[65]), .s(stg1_s7[66]), .c(stg1_c7[66]), .co(stg1_co7[66]));
counter_5to3 u_a17_67(.i0(pp25_w[65]), .i1(pp26_w[65]), .i2(pp27_w[63]), .i3(pp28_w[61]), .ci(stg1_co7[66]), .s(stg1_s7[67]), .c(stg1_c7[67]), .co(stg1_co7[67]));
counter_5to3 u_a17_68(.i0(pp25_w[65]), .i1(pp26_w[65]), .i2(pp27_w[64]), .i3(pp28_w[62]), .ci(stg1_co7[67]), .s(stg1_s7[68]), .c(stg1_c7[68]), .co(stg1_co7[68]));
counter_5to3 u_a17_69(.i0(pp25_w[65]), .i1(pp26_w[65]), .i2(pp27_w[65]), .i3(pp28_w[63]), .ci(stg1_co7[68]), .s(stg1_s7[69]), .c(stg1_c7[69]), .co(stg1_co7[69]));
counter_5to3 u_a17_70(.i0(pp25_w[65]), .i1(pp26_w[65]), .i2(pp27_w[65]), .i3(pp28_w[64]), .ci(stg1_co7[69]), .s(stg1_s7[70]), .c(stg1_c7[70]), .co(stg1_co7[70]));
counter_5to3 u_al7_71(.i0(pp25_w[65]), .i1(pp26_w[65]), .i2(pp27_w[65]), .i3(pp28_w[65]), .ci(stg1_co7[70]), .s(stg1_s7[71]), .c(stg1_c7[71]), .co(stg1_co7[71]));
counter_5to3 u_al7_72(.i0(pp25_w[65]), .i1(pp26_w[65]), .i2(pp27_w[65]), .i3(pp28_w[65]), .ci(stg1_co7[71]), .s(stg1_s7[72]), .c(stg1_c7[72]), .co(stg1_co7[72]));

// =========================== first stage 8th group ============================================================================================================
counter_5to3 u_a18_0 (.i0(pp29_w[0 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(1'b0        ), .s(stg1_s8[0 ]), .c(stg1_c8[0 ]), .co(stg1_co8[0 ]));
counter_5to3 u_a18_1 (.i0(pp29_w[1 ]), .i1(1'b0      ), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co8[0 ]), .s(stg1_s8[1 ]), .c(stg1_c8[1 ]), .co(stg1_co8[1 ]));
counter_5to3 u_a18_2 (.i0(pp29_w[2 ]), .i1(pp30_w[0 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co8[1 ]), .s(stg1_s8[2 ]), .c(stg1_c8[2 ]), .co(stg1_co8[2 ]));
counter_5to3 u_a18_3 (.i0(pp29_w[3 ]), .i1(pp30_w[1 ]), .i2(1'b0      ), .i3(1'b0      ), .ci(stg1_co8[2 ]), .s(stg1_s8[3 ]), .c(stg1_c8[3 ]), .co(stg1_co8[3 ]));
counter_5to3 u_a18_4 (.i0(pp29_w[4 ]), .i1(pp30_w[2 ]), .i2(pp31_w[0 ]), .i3(1'b0      ), .ci(stg1_co8[3 ]), .s(stg1_s8[4 ]), .c(stg1_c8[4 ]), .co(stg1_co8[4 ]));
counter_5to3 u_a18_5 (.i0(pp29_w[5 ]), .i1(pp30_w[3 ]), .i2(pp31_w[1 ]), .i3(1'b0      ), .ci(stg1_co8[4 ]), .s(stg1_s8[5 ]), .c(stg1_c8[5 ]), .co(stg1_co8[5 ]));
counter_5to3 u_a18_6 (.i0(pp29_w[6 ]), .i1(pp30_w[4 ]), .i2(pp31_w[2 ]), .i3(pp32_w[0 ]), .ci(stg1_co8[5 ]), .s(stg1_s8[6 ]), .c(stg1_c8[6 ]), .co(stg1_co8[6 ]));
counter_5to3 u_a18_7 (.i0(pp29_w[7 ]), .i1(pp30_w[5 ]), .i2(pp31_w[3 ]), .i3(pp32_w[1 ]), .ci(stg1_co8[6 ]), .s(stg1_s8[7 ]), .c(stg1_c8[7 ]), .co(stg1_co8[7 ]));
counter_5to3 u_a18_8 (.i0(pp29_w[8 ]), .i1(pp30_w[6 ]), .i2(pp31_w[4 ]), .i3(pp32_w[2 ]), .ci(stg1_co8[7 ]), .s(stg1_s8[8 ]), .c(stg1_c8[8 ]), .co(stg1_co8[8 ]));
counter_5to3 u_a18_9 (.i0(pp29_w[9 ]), .i1(pp30_w[7 ]), .i2(pp31_w[5 ]), .i3(pp32_w[3 ]), .ci(stg1_co8[8 ]), .s(stg1_s8[9 ]), .c(stg1_c8[9 ]), .co(stg1_co8[9 ]));
counter_5to3 u_a18_10(.i0(pp29_w[10]), .i1(pp30_w[8 ]), .i2(pp31_w[6 ]), .i3(pp32_w[4 ]), .ci(stg1_co8[9 ]), .s(stg1_s8[10]), .c(stg1_c8[10]), .co(stg1_co8[10]));
counter_5to3 u_a18_11(.i0(pp29_w[11]), .i1(pp30_w[9 ]), .i2(pp31_w[7 ]), .i3(pp32_w[5 ]), .ci(stg1_co8[10]), .s(stg1_s8[11]), .c(stg1_c8[11]), .co(stg1_co8[11]));
counter_5to3 u_a18_12(.i0(pp29_w[12]), .i1(pp30_w[10]), .i2(pp31_w[8 ]), .i3(pp32_w[6 ]), .ci(stg1_co8[11]), .s(stg1_s8[12]), .c(stg1_c8[12]), .co(stg1_co8[12]));
counter_5to3 u_a18_13(.i0(pp29_w[13]), .i1(pp30_w[11]), .i2(pp31_w[9 ]), .i3(pp32_w[7 ]), .ci(stg1_co8[12]), .s(stg1_s8[13]), .c(stg1_c8[13]), .co(stg1_co8[13]));
counter_5to3 u_a18_14(.i0(pp29_w[14]), .i1(pp30_w[12]), .i2(pp31_w[10]), .i3(pp32_w[8 ]), .ci(stg1_co8[13]), .s(stg1_s8[14]), .c(stg1_c8[14]), .co(stg1_co8[14]));
counter_5to3 u_a18_15(.i0(pp29_w[15]), .i1(pp30_w[13]), .i2(pp31_w[11]), .i3(pp32_w[9 ]), .ci(stg1_co8[14]), .s(stg1_s8[15]), .c(stg1_c8[15]), .co(stg1_co8[15]));
counter_5to3 u_a18_16(.i0(pp29_w[16]), .i1(pp30_w[14]), .i2(pp31_w[12]), .i3(pp32_w[10]), .ci(stg1_co8[15]), .s(stg1_s8[16]), .c(stg1_c8[16]), .co(stg1_co8[16]));
counter_5to3 u_a18_17(.i0(pp29_w[17]), .i1(pp30_w[15]), .i2(pp31_w[13]), .i3(pp32_w[11]), .ci(stg1_co8[16]), .s(stg1_s8[17]), .c(stg1_c8[17]), .co(stg1_co8[17]));
counter_5to3 u_a18_18(.i0(pp29_w[18]), .i1(pp30_w[16]), .i2(pp31_w[14]), .i3(pp32_w[12]), .ci(stg1_co8[17]), .s(stg1_s8[18]), .c(stg1_c8[18]), .co(stg1_co8[18]));
counter_5to3 u_a18_19(.i0(pp29_w[19]), .i1(pp30_w[17]), .i2(pp31_w[15]), .i3(pp32_w[13]), .ci(stg1_co8[18]), .s(stg1_s8[19]), .c(stg1_c8[19]), .co(stg1_co8[19]));
counter_5to3 u_a18_20(.i0(pp29_w[20]), .i1(pp30_w[18]), .i2(pp31_w[16]), .i3(pp32_w[14]), .ci(stg1_co8[19]), .s(stg1_s8[20]), .c(stg1_c8[20]), .co(stg1_co8[20]));
counter_5to3 u_a18_21(.i0(pp29_w[21]), .i1(pp30_w[19]), .i2(pp31_w[17]), .i3(pp32_w[15]), .ci(stg1_co8[20]), .s(stg1_s8[21]), .c(stg1_c8[21]), .co(stg1_co8[21]));
counter_5to3 u_a18_22(.i0(pp29_w[22]), .i1(pp30_w[20]), .i2(pp31_w[18]), .i3(pp32_w[16]), .ci(stg1_co8[21]), .s(stg1_s8[22]), .c(stg1_c8[22]), .co(stg1_co8[22]));
counter_5to3 u_a18_23(.i0(pp29_w[23]), .i1(pp30_w[21]), .i2(pp31_w[19]), .i3(pp32_w[17]), .ci(stg1_co8[22]), .s(stg1_s8[23]), .c(stg1_c8[23]), .co(stg1_co8[23]));
counter_5to3 u_a18_24(.i0(pp29_w[24]), .i1(pp30_w[22]), .i2(pp31_w[20]), .i3(pp32_w[18]), .ci(stg1_co8[23]), .s(stg1_s8[24]), .c(stg1_c8[24]), .co(stg1_co8[24]));
counter_5to3 u_a18_25(.i0(pp29_w[25]), .i1(pp30_w[23]), .i2(pp31_w[21]), .i3(pp32_w[19]), .ci(stg1_co8[24]), .s(stg1_s8[25]), .c(stg1_c8[25]), .co(stg1_co8[25]));
counter_5to3 u_a18_26(.i0(pp29_w[26]), .i1(pp30_w[24]), .i2(pp31_w[22]), .i3(pp32_w[20]), .ci(stg1_co8[25]), .s(stg1_s8[26]), .c(stg1_c8[26]), .co(stg1_co8[26]));
counter_5to3 u_a18_27(.i0(pp29_w[27]), .i1(pp30_w[25]), .i2(pp31_w[23]), .i3(pp32_w[21]), .ci(stg1_co8[26]), .s(stg1_s8[27]), .c(stg1_c8[27]), .co(stg1_co8[27]));
counter_5to3 u_a18_28(.i0(pp29_w[28]), .i1(pp30_w[26]), .i2(pp31_w[24]), .i3(pp32_w[22]), .ci(stg1_co8[27]), .s(stg1_s8[28]), .c(stg1_c8[28]), .co(stg1_co8[28]));
counter_5to3 u_a18_29(.i0(pp29_w[29]), .i1(pp30_w[27]), .i2(pp31_w[25]), .i3(pp32_w[23]), .ci(stg1_co8[28]), .s(stg1_s8[29]), .c(stg1_c8[29]), .co(stg1_co8[29]));
counter_5to3 u_a18_30(.i0(pp29_w[30]), .i1(pp30_w[28]), .i2(pp31_w[26]), .i3(pp32_w[24]), .ci(stg1_co8[29]), .s(stg1_s8[30]), .c(stg1_c8[30]), .co(stg1_co8[30]));
counter_5to3 u_a18_31(.i0(pp29_w[31]), .i1(pp30_w[29]), .i2(pp31_w[27]), .i3(pp32_w[25]), .ci(stg1_co8[30]), .s(stg1_s8[31]), .c(stg1_c8[31]), .co(stg1_co8[31]));
counter_5to3 u_a18_32(.i0(pp29_w[32]), .i1(pp30_w[30]), .i2(pp31_w[28]), .i3(pp32_w[26]), .ci(stg1_co8[31]), .s(stg1_s8[32]), .c(stg1_c8[32]), .co(stg1_co8[32]));
counter_5to3 u_a18_33(.i0(pp29_w[33]), .i1(pp30_w[31]), .i2(pp31_w[29]), .i3(pp32_w[27]), .ci(stg1_co8[32]), .s(stg1_s8[33]), .c(stg1_c8[33]), .co(stg1_co8[33]));
counter_5to3 u_a18_34(.i0(pp29_w[34]), .i1(pp30_w[32]), .i2(pp31_w[30]), .i3(pp32_w[28]), .ci(stg1_co8[33]), .s(stg1_s8[34]), .c(stg1_c8[34]), .co(stg1_co8[34]));
counter_5to3 u_a18_35(.i0(pp29_w[35]), .i1(pp30_w[33]), .i2(pp31_w[31]), .i3(pp32_w[29]), .ci(stg1_co8[34]), .s(stg1_s8[35]), .c(stg1_c8[35]), .co(stg1_co8[35]));
counter_5to3 u_a18_36(.i0(pp29_w[36]), .i1(pp30_w[34]), .i2(pp31_w[32]), .i3(pp32_w[30]), .ci(stg1_co8[35]), .s(stg1_s8[36]), .c(stg1_c8[36]), .co(stg1_co8[36]));
counter_5to3 u_a18_37(.i0(pp29_w[37]), .i1(pp30_w[35]), .i2(pp31_w[33]), .i3(pp32_w[31]), .ci(stg1_co8[36]), .s(stg1_s8[37]), .c(stg1_c8[37]), .co(stg1_co8[37]));
counter_5to3 u_a18_38(.i0(pp29_w[38]), .i1(pp30_w[36]), .i2(pp31_w[34]), .i3(pp32_w[32]), .ci(stg1_co8[37]), .s(stg1_s8[38]), .c(stg1_c8[38]), .co(stg1_co8[38]));
counter_5to3 u_a18_39(.i0(pp29_w[39]), .i1(pp30_w[37]), .i2(pp31_w[35]), .i3(pp32_w[33]), .ci(stg1_co8[38]), .s(stg1_s8[39]), .c(stg1_c8[39]), .co(stg1_co8[39]));
counter_5to3 u_a18_40(.i0(pp29_w[40]), .i1(pp30_w[38]), .i2(pp31_w[36]), .i3(pp32_w[34]), .ci(stg1_co8[39]), .s(stg1_s8[40]), .c(stg1_c8[40]), .co(stg1_co8[40]));
counter_5to3 u_a18_41(.i0(pp29_w[41]), .i1(pp30_w[39]), .i2(pp31_w[37]), .i3(pp32_w[35]), .ci(stg1_co8[40]), .s(stg1_s8[41]), .c(stg1_c8[41]), .co(stg1_co8[41]));
counter_5to3 u_a18_42(.i0(pp29_w[42]), .i1(pp30_w[40]), .i2(pp31_w[38]), .i3(pp32_w[36]), .ci(stg1_co8[41]), .s(stg1_s8[42]), .c(stg1_c8[42]), .co(stg1_co8[42]));
counter_5to3 u_a18_43(.i0(pp29_w[43]), .i1(pp30_w[41]), .i2(pp31_w[39]), .i3(pp32_w[37]), .ci(stg1_co8[42]), .s(stg1_s8[43]), .c(stg1_c8[43]), .co(stg1_co8[43]));
counter_5to3 u_a18_44(.i0(pp29_w[44]), .i1(pp30_w[42]), .i2(pp31_w[40]), .i3(pp32_w[38]), .ci(stg1_co8[43]), .s(stg1_s8[44]), .c(stg1_c8[44]), .co(stg1_co8[44]));
counter_5to3 u_a18_45(.i0(pp29_w[45]), .i1(pp30_w[43]), .i2(pp31_w[41]), .i3(pp32_w[39]), .ci(stg1_co8[44]), .s(stg1_s8[45]), .c(stg1_c8[45]), .co(stg1_co8[45]));
counter_5to3 u_a18_46(.i0(pp29_w[46]), .i1(pp30_w[44]), .i2(pp31_w[42]), .i3(pp32_w[40]), .ci(stg1_co8[45]), .s(stg1_s8[46]), .c(stg1_c8[46]), .co(stg1_co8[46]));
counter_5to3 u_a18_47(.i0(pp29_w[47]), .i1(pp30_w[45]), .i2(pp31_w[43]), .i3(pp32_w[41]), .ci(stg1_co8[46]), .s(stg1_s8[47]), .c(stg1_c8[47]), .co(stg1_co8[47]));
counter_5to3 u_a18_48(.i0(pp29_w[48]), .i1(pp30_w[46]), .i2(pp31_w[44]), .i3(pp32_w[42]), .ci(stg1_co8[47]), .s(stg1_s8[48]), .c(stg1_c8[48]), .co(stg1_co8[48]));
counter_5to3 u_a18_49(.i0(pp29_w[49]), .i1(pp30_w[47]), .i2(pp31_w[45]), .i3(pp32_w[43]), .ci(stg1_co8[48]), .s(stg1_s8[49]), .c(stg1_c8[49]), .co(stg1_co8[49]));
counter_5to3 u_a18_50(.i0(pp29_w[50]), .i1(pp30_w[48]), .i2(pp31_w[46]), .i3(pp32_w[44]), .ci(stg1_co8[49]), .s(stg1_s8[50]), .c(stg1_c8[50]), .co(stg1_co8[50]));
counter_5to3 u_a18_51(.i0(pp29_w[51]), .i1(pp30_w[49]), .i2(pp31_w[47]), .i3(pp32_w[45]), .ci(stg1_co8[50]), .s(stg1_s8[51]), .c(stg1_c8[51]), .co(stg1_co8[51]));
counter_5to3 u_a18_52(.i0(pp29_w[52]), .i1(pp30_w[50]), .i2(pp31_w[48]), .i3(pp32_w[46]), .ci(stg1_co8[51]), .s(stg1_s8[52]), .c(stg1_c8[52]), .co(stg1_co8[52]));
counter_5to3 u_a18_53(.i0(pp29_w[53]), .i1(pp30_w[51]), .i2(pp31_w[49]), .i3(pp32_w[47]), .ci(stg1_co8[52]), .s(stg1_s8[53]), .c(stg1_c8[53]), .co(stg1_co8[53]));
counter_5to3 u_a18_54(.i0(pp29_w[54]), .i1(pp30_w[52]), .i2(pp31_w[50]), .i3(pp32_w[48]), .ci(stg1_co8[53]), .s(stg1_s8[54]), .c(stg1_c8[54]), .co(stg1_co8[54]));
counter_5to3 u_a18_55(.i0(pp29_w[55]), .i1(pp30_w[53]), .i2(pp31_w[51]), .i3(pp32_w[49]), .ci(stg1_co8[54]), .s(stg1_s8[55]), .c(stg1_c8[55]), .co(stg1_co8[55]));
counter_5to3 u_a18_56(.i0(pp29_w[56]), .i1(pp30_w[54]), .i2(pp31_w[52]), .i3(pp32_w[50]), .ci(stg1_co8[55]), .s(stg1_s8[56]), .c(stg1_c8[56]), .co(stg1_co8[56]));
counter_5to3 u_a18_57(.i0(pp29_w[57]), .i1(pp30_w[55]), .i2(pp31_w[53]), .i3(pp32_w[51]), .ci(stg1_co8[56]), .s(stg1_s8[57]), .c(stg1_c8[57]), .co(stg1_co8[57]));
counter_5to3 u_a18_58(.i0(pp29_w[58]), .i1(pp30_w[56]), .i2(pp31_w[54]), .i3(pp32_w[52]), .ci(stg1_co8[57]), .s(stg1_s8[58]), .c(stg1_c8[58]), .co(stg1_co8[58]));
counter_5to3 u_a18_59(.i0(pp29_w[59]), .i1(pp30_w[57]), .i2(pp31_w[55]), .i3(pp32_w[53]), .ci(stg1_co8[58]), .s(stg1_s8[59]), .c(stg1_c8[59]), .co(stg1_co8[59]));
counter_5to3 u_a18_60(.i0(pp29_w[60]), .i1(pp30_w[58]), .i2(pp31_w[56]), .i3(pp32_w[54]), .ci(stg1_co8[59]), .s(stg1_s8[60]), .c(stg1_c8[60]), .co(stg1_co8[60]));
counter_5to3 u_a18_61(.i0(pp29_w[61]), .i1(pp30_w[59]), .i2(pp31_w[57]), .i3(pp32_w[55]), .ci(stg1_co8[60]), .s(stg1_s8[61]), .c(stg1_c8[61]), .co(stg1_co8[61]));
counter_5to3 u_a18_62(.i0(pp29_w[62]), .i1(pp30_w[60]), .i2(pp31_w[58]), .i3(pp32_w[56]), .ci(stg1_co8[61]), .s(stg1_s8[62]), .c(stg1_c8[62]), .co(stg1_co8[62]));
counter_5to3 u_a18_63(.i0(pp29_w[63]), .i1(pp30_w[61]), .i2(pp31_w[59]), .i3(pp32_w[57]), .ci(stg1_co8[62]), .s(stg1_s8[63]), .c(stg1_c8[63]), .co(stg1_co8[63]));
counter_5to3 u_a18_64(.i0(pp29_w[64]), .i1(pp30_w[62]), .i2(pp31_w[60]), .i3(pp32_w[58]), .ci(stg1_co8[63]), .s(stg1_s8[64]), .c(stg1_c8[64]), .co(stg1_co8[64]));
counter_5to3 u_a18_65(.i0(pp29_w[65]), .i1(pp30_w[63]), .i2(pp31_w[61]), .i3(pp32_w[59]), .ci(stg1_co8[64]), .s(stg1_s8[65]), .c(stg1_c8[65]), .co(stg1_co8[65]));
counter_5to3 u_a18_66(.i0(pp29_w[65]), .i1(pp30_w[64]), .i2(pp31_w[62]), .i3(pp32_w[60]), .ci(stg1_co8[65]), .s(stg1_s8[66]), .c(stg1_c8[66]), .co(stg1_co8[66]));
counter_5to3 u_a18_67(.i0(pp29_w[65]), .i1(pp30_w[65]), .i2(pp31_w[63]), .i3(pp32_w[61]), .ci(stg1_co8[66]), .s(stg1_s8[67]), .c(stg1_c8[67]), .co(stg1_co8[67]));
counter_5to3 u_a18_68(.i0(pp29_w[65]), .i1(pp30_w[65]), .i2(pp31_w[64]), .i3(pp32_w[62]), .ci(stg1_co8[67]), .s(stg1_s8[68]), .c(stg1_c8[68]), .co(stg1_co8[68]));
counter_5to3 u_a18_69(.i0(pp29_w[65]), .i1(pp30_w[65]), .i2(pp31_w[65]), .i3(pp32_w[63]), .ci(stg1_co8[68]), .s(stg1_s8[69]), .c(stg1_c8[69]), .co(stg1_co8[69]));
counter_5to3 u_a18_70(.i0(pp29_w[65]), .i1(pp30_w[65]), .i2(pp31_w[65]), .i3(pp32_w[64]), .ci(stg1_co8[69]), .s(stg1_s8[70]), .c(stg1_c8[70]), .co(stg1_co8[70]));
counter_5to3 u_al8_71(.i0(pp29_w[65]), .i1(pp30_w[65]), .i2(pp31_w[65]), .i3(pp32_w[65]), .ci(stg1_co8[70]), .s(stg1_s8[71]), .c(stg1_c8[71]), .co(stg1_co8[71]));

//================ second stage ================
wire [72:0] stg1_s1_w, stg1_c1_w;
wire [72:0] stg1_s2_w, stg1_c2_w;
wire [72:0] stg1_s3_w, stg1_c3_w;
wire [72:0] stg1_s4_w, stg1_c4_w;
wire [72:0] stg1_s5_w, stg1_c5_w;
wire [72:0] stg1_s6_w, stg1_c6_w;
wire [72:0] stg1_s7_w, stg1_c7_w;
wire [71:0] stg1_s8_w, stg1_c8_w;
wire [65:0] pp33_w1;

// ============= pipeline ===============
reg [72:0] stg1_s1_ff, stg1_c1_ff;
reg [72:0] stg1_s2_ff, stg1_c2_ff;
reg [72:0] stg1_s3_ff, stg1_c3_ff;
reg [72:0] stg1_s4_ff, stg1_c4_ff;
reg [72:0] stg1_s5_ff, stg1_c5_ff;
reg [72:0] stg1_s6_ff, stg1_c6_ff;
reg [72:0] stg1_s7_ff, stg1_c7_ff;
reg [71:0] stg1_s8_ff, stg1_c8_ff;
reg [65:0] pp33_f1;

always @(posedge clk or negedge rstn)begin
    if (!rstn)begin
        stg1_s1_ff <= 73'b0;
        stg1_c1_ff <= 73'b0;
        stg1_s2_ff <= 73'b0;
        stg1_c2_ff <= 73'b0;
        stg1_s3_ff <= 73'b0;
        stg1_c3_ff <= 73'b0;
        stg1_s4_ff <= 73'b0;
        stg1_c4_ff <= 73'b0;
        stg1_s5_ff <= 73'b0;
        stg1_c5_ff <= 73'b0;
        stg1_s6_ff <= 73'b0;
        stg1_c6_ff <= 73'b0;
        stg1_s7_ff <= 73'b0;
        stg1_c7_ff <= 73'b0;
        stg1_s8_ff <= 72'b0;
        stg1_c8_ff <= 72'b0;
        pp33_f1    <= 66'b0;
    end
    else begin
        stg1_s1_ff   <= stg1_s1;
        stg1_c1_ff   <= stg1_c1;
        stg1_s2_ff   <= stg1_s2;
        stg1_c2_ff   <= stg1_c2;
        stg1_s3_ff   <= stg1_s3;
        stg1_c3_ff   <= stg1_c3;
        stg1_s4_ff   <= stg1_s4;
        stg1_c4_ff   <= stg1_c4;
        stg1_s5_ff   <= stg1_s5;
        stg1_c5_ff   <= stg1_c5;
        stg1_s6_ff   <= stg1_s6;
        stg1_c6_ff   <= stg1_c6;
        stg1_s7_ff   <= stg1_s7;
        stg1_c7_ff   <= stg1_c7;
        stg1_s8_ff   <= stg1_s8;
        stg1_c8_ff   <= stg1_c8;
        pp33_f1      <= pp33_w;
    end
end

assign stg1_s1_w   = stg1_s1_ff;
assign stg1_c1_w   = stg1_c1_ff;
assign stg1_s2_w   = stg1_s2_ff;
assign stg1_c2_w   = stg1_c2_ff;
assign stg1_s3_w   = stg1_s3_ff;
assign stg1_c3_w   = stg1_c3_ff;
assign stg1_s4_w   = stg1_s4_ff;
assign stg1_c4_w   = stg1_c4_ff;
assign stg1_s5_w   = stg1_s5_ff;
assign stg1_c5_w   = stg1_c5_ff;
assign stg1_s6_w   = stg1_s6_ff;
assign stg1_c6_w   = stg1_c6_ff;
assign stg1_s7_w   = stg1_s7_ff;
assign stg1_c7_w   = stg1_c7_ff;
assign stg1_s8_w   = stg1_s8_ff;
assign stg1_c8_w   = stg1_c8_ff;
assign pp33_w1     = pp33_f1   ;

wire [82:0] stg2_s1, stg2_c1, stg2_co1;
wire [82:0] stg2_s2, stg2_c2, stg2_co2;
wire [82:0] stg2_s3, stg2_c3, stg2_co3;
wire [79:0] stg2_s4, stg2_c4, stg2_co4;

// =========================== second stage 1st group ============================================================================================================
counter_5to3 u_a21_0 (.i0(stg1_s1_w[0 ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0         ), .ci(1'b0        ), .s(stg2_s1[0 ]), .c(stg2_c1[0 ]), .co(stg2_co1[0 ]));
counter_5to3 u_a21_1 (.i0(stg1_s1_w[1 ]), .i1(stg1_c1_w[0 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[0 ]), .s(stg2_s1[1 ]), .c(stg2_c1[1 ]), .co(stg2_co1[1 ]));
counter_5to3 u_a21_2 (.i0(stg1_s1_w[2 ]), .i1(stg1_c1_w[1 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[1 ]), .s(stg2_s1[2 ]), .c(stg2_c1[2 ]), .co(stg2_co1[2 ]));
counter_5to3 u_a21_3 (.i0(stg1_s1_w[3 ]), .i1(stg1_c1_w[2 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[2 ]), .s(stg2_s1[3 ]), .c(stg2_c1[3 ]), .co(stg2_co1[3 ]));
counter_5to3 u_a21_4 (.i0(stg1_s1_w[4 ]), .i1(stg1_c1_w[3 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[3 ]), .s(stg2_s1[4 ]), .c(stg2_c1[4 ]), .co(stg2_co1[4 ]));
counter_5to3 u_a21_5 (.i0(stg1_s1_w[5 ]), .i1(stg1_c1_w[4 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[4 ]), .s(stg2_s1[5 ]), .c(stg2_c1[5 ]), .co(stg2_co1[5 ]));
counter_5to3 u_a21_6 (.i0(stg1_s1_w[6 ]), .i1(stg1_c1_w[5 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[5 ]), .s(stg2_s1[6 ]), .c(stg2_c1[6 ]), .co(stg2_co1[6 ]));
counter_5to3 u_a21_7 (.i0(stg1_s1_w[7 ]), .i1(stg1_c1_w[6 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co1[6 ]), .s(stg2_s1[7 ]), .c(stg2_c1[7 ]), .co(stg2_co1[7 ]));
counter_5to3 u_a21_8 (.i0(stg1_s1_w[8 ]), .i1(stg1_c1_w[7 ]), .i2(stg1_s2_w[0 ]), .i3(1'b0         ), .ci(stg2_co1[7 ]), .s(stg2_s1[8 ]), .c(stg2_c1[8 ]), .co(stg2_co1[8 ]));
counter_5to3 u_a21_9 (.i0(stg1_s1_w[9 ]), .i1(stg1_c1_w[8 ]), .i2(stg1_s2_w[1 ]), .i3(stg1_c2_w[0 ]), .ci(stg2_co1[8 ]), .s(stg2_s1[9 ]), .c(stg2_c1[9 ]), .co(stg2_co1[9 ]));
counter_5to3 u_a21_10(.i0(stg1_s1_w[10]), .i1(stg1_c1_w[9 ]), .i2(stg1_s2_w[2 ]), .i3(stg1_c2_w[1 ]), .ci(stg2_co1[9 ]), .s(stg2_s1[10]), .c(stg2_c1[10]), .co(stg2_co1[10]));
counter_5to3 u_a21_11(.i0(stg1_s1_w[11]), .i1(stg1_c1_w[10]), .i2(stg1_s2_w[3 ]), .i3(stg1_c2_w[2 ]), .ci(stg2_co1[10]), .s(stg2_s1[11]), .c(stg2_c1[11]), .co(stg2_co1[11]));
counter_5to3 u_a21_12(.i0(stg1_s1_w[12]), .i1(stg1_c1_w[11]), .i2(stg1_s2_w[4 ]), .i3(stg1_c2_w[3 ]), .ci(stg2_co1[11]), .s(stg2_s1[12]), .c(stg2_c1[12]), .co(stg2_co1[12]));
counter_5to3 u_a21_13(.i0(stg1_s1_w[13]), .i1(stg1_c1_w[12]), .i2(stg1_s2_w[5 ]), .i3(stg1_c2_w[4 ]), .ci(stg2_co1[12]), .s(stg2_s1[13]), .c(stg2_c1[13]), .co(stg2_co1[13]));
counter_5to3 u_a21_14(.i0(stg1_s1_w[14]), .i1(stg1_c1_w[13]), .i2(stg1_s2_w[6 ]), .i3(stg1_c2_w[5 ]), .ci(stg2_co1[13]), .s(stg2_s1[14]), .c(stg2_c1[14]), .co(stg2_co1[14]));
counter_5to3 u_a21_15(.i0(stg1_s1_w[15]), .i1(stg1_c1_w[14]), .i2(stg1_s2_w[7 ]), .i3(stg1_c2_w[6 ]), .ci(stg2_co1[14]), .s(stg2_s1[15]), .c(stg2_c1[15]), .co(stg2_co1[15]));
counter_5to3 u_a21_16(.i0(stg1_s1_w[16]), .i1(stg1_c1_w[15]), .i2(stg1_s2_w[8 ]), .i3(stg1_c2_w[7 ]), .ci(stg2_co1[15]), .s(stg2_s1[16]), .c(stg2_c1[16]), .co(stg2_co1[16]));
counter_5to3 u_a21_17(.i0(stg1_s1_w[17]), .i1(stg1_c1_w[16]), .i2(stg1_s2_w[9 ]), .i3(stg1_c2_w[8 ]), .ci(stg2_co1[16]), .s(stg2_s1[17]), .c(stg2_c1[17]), .co(stg2_co1[17]));
counter_5to3 u_a21_18(.i0(stg1_s1_w[18]), .i1(stg1_c1_w[17]), .i2(stg1_s2_w[10]), .i3(stg1_c2_w[9 ]), .ci(stg2_co1[17]), .s(stg2_s1[18]), .c(stg2_c1[18]), .co(stg2_co1[18]));
counter_5to3 u_a21_19(.i0(stg1_s1_w[19]), .i1(stg1_c1_w[18]), .i2(stg1_s2_w[11]), .i3(stg1_c2_w[10]), .ci(stg2_co1[18]), .s(stg2_s1[19]), .c(stg2_c1[19]), .co(stg2_co1[19]));
counter_5to3 u_a21_20(.i0(stg1_s1_w[20]), .i1(stg1_c1_w[19]), .i2(stg1_s2_w[12]), .i3(stg1_c2_w[11]), .ci(stg2_co1[19]), .s(stg2_s1[20]), .c(stg2_c1[20]), .co(stg2_co1[20]));
counter_5to3 u_a21_21(.i0(stg1_s1_w[21]), .i1(stg1_c1_w[20]), .i2(stg1_s2_w[13]), .i3(stg1_c2_w[12]), .ci(stg2_co1[20]), .s(stg2_s1[21]), .c(stg2_c1[21]), .co(stg2_co1[21]));
counter_5to3 u_a21_22(.i0(stg1_s1_w[22]), .i1(stg1_c1_w[21]), .i2(stg1_s2_w[14]), .i3(stg1_c2_w[13]), .ci(stg2_co1[21]), .s(stg2_s1[22]), .c(stg2_c1[22]), .co(stg2_co1[22]));
counter_5to3 u_a21_23(.i0(stg1_s1_w[23]), .i1(stg1_c1_w[22]), .i2(stg1_s2_w[15]), .i3(stg1_c2_w[14]), .ci(stg2_co1[22]), .s(stg2_s1[23]), .c(stg2_c1[23]), .co(stg2_co1[23]));
counter_5to3 u_a21_24(.i0(stg1_s1_w[24]), .i1(stg1_c1_w[23]), .i2(stg1_s2_w[16]), .i3(stg1_c2_w[15]), .ci(stg2_co1[23]), .s(stg2_s1[24]), .c(stg2_c1[24]), .co(stg2_co1[24]));
counter_5to3 u_a21_25(.i0(stg1_s1_w[25]), .i1(stg1_c1_w[24]), .i2(stg1_s2_w[17]), .i3(stg1_c2_w[16]), .ci(stg2_co1[24]), .s(stg2_s1[25]), .c(stg2_c1[25]), .co(stg2_co1[25]));
counter_5to3 u_a21_26(.i0(stg1_s1_w[26]), .i1(stg1_c1_w[25]), .i2(stg1_s2_w[18]), .i3(stg1_c2_w[17]), .ci(stg2_co1[25]), .s(stg2_s1[26]), .c(stg2_c1[26]), .co(stg2_co1[26]));
counter_5to3 u_a21_27(.i0(stg1_s1_w[27]), .i1(stg1_c1_w[26]), .i2(stg1_s2_w[19]), .i3(stg1_c2_w[18]), .ci(stg2_co1[26]), .s(stg2_s1[27]), .c(stg2_c1[27]), .co(stg2_co1[27]));
counter_5to3 u_a21_28(.i0(stg1_s1_w[28]), .i1(stg1_c1_w[27]), .i2(stg1_s2_w[20]), .i3(stg1_c2_w[19]), .ci(stg2_co1[27]), .s(stg2_s1[28]), .c(stg2_c1[28]), .co(stg2_co1[28]));
counter_5to3 u_a21_29(.i0(stg1_s1_w[29]), .i1(stg1_c1_w[28]), .i2(stg1_s2_w[21]), .i3(stg1_c2_w[20]), .ci(stg2_co1[28]), .s(stg2_s1[29]), .c(stg2_c1[29]), .co(stg2_co1[29]));
counter_5to3 u_a21_30(.i0(stg1_s1_w[30]), .i1(stg1_c1_w[29]), .i2(stg1_s2_w[22]), .i3(stg1_c2_w[21]), .ci(stg2_co1[29]), .s(stg2_s1[30]), .c(stg2_c1[30]), .co(stg2_co1[30]));
counter_5to3 u_a21_31(.i0(stg1_s1_w[31]), .i1(stg1_c1_w[30]), .i2(stg1_s2_w[23]), .i3(stg1_c2_w[22]), .ci(stg2_co1[30]), .s(stg2_s1[31]), .c(stg2_c1[31]), .co(stg2_co1[31]));
counter_5to3 u_a21_32(.i0(stg1_s1_w[32]), .i1(stg1_c1_w[31]), .i2(stg1_s2_w[24]), .i3(stg1_c2_w[23]), .ci(stg2_co1[31]), .s(stg2_s1[32]), .c(stg2_c1[32]), .co(stg2_co1[32]));
counter_5to3 u_a21_33(.i0(stg1_s1_w[33]), .i1(stg1_c1_w[32]), .i2(stg1_s2_w[25]), .i3(stg1_c2_w[24]), .ci(stg2_co1[32]), .s(stg2_s1[33]), .c(stg2_c1[33]), .co(stg2_co1[33]));
counter_5to3 u_a21_34(.i0(stg1_s1_w[34]), .i1(stg1_c1_w[33]), .i2(stg1_s2_w[26]), .i3(stg1_c2_w[25]), .ci(stg2_co1[33]), .s(stg2_s1[34]), .c(stg2_c1[34]), .co(stg2_co1[34]));
counter_5to3 u_a21_35(.i0(stg1_s1_w[35]), .i1(stg1_c1_w[34]), .i2(stg1_s2_w[27]), .i3(stg1_c2_w[26]), .ci(stg2_co1[34]), .s(stg2_s1[35]), .c(stg2_c1[35]), .co(stg2_co1[35]));
counter_5to3 u_a21_36(.i0(stg1_s1_w[36]), .i1(stg1_c1_w[35]), .i2(stg1_s2_w[28]), .i3(stg1_c2_w[27]), .ci(stg2_co1[35]), .s(stg2_s1[36]), .c(stg2_c1[36]), .co(stg2_co1[36]));
counter_5to3 u_a21_37(.i0(stg1_s1_w[37]), .i1(stg1_c1_w[36]), .i2(stg1_s2_w[29]), .i3(stg1_c2_w[28]), .ci(stg2_co1[36]), .s(stg2_s1[37]), .c(stg2_c1[37]), .co(stg2_co1[37]));
counter_5to3 u_a21_38(.i0(stg1_s1_w[38]), .i1(stg1_c1_w[37]), .i2(stg1_s2_w[30]), .i3(stg1_c2_w[29]), .ci(stg2_co1[37]), .s(stg2_s1[38]), .c(stg2_c1[38]), .co(stg2_co1[38]));
counter_5to3 u_a21_39(.i0(stg1_s1_w[39]), .i1(stg1_c1_w[38]), .i2(stg1_s2_w[31]), .i3(stg1_c2_w[30]), .ci(stg2_co1[38]), .s(stg2_s1[39]), .c(stg2_c1[39]), .co(stg2_co1[39]));
counter_5to3 u_a21_40(.i0(stg1_s1_w[40]), .i1(stg1_c1_w[39]), .i2(stg1_s2_w[32]), .i3(stg1_c2_w[31]), .ci(stg2_co1[39]), .s(stg2_s1[40]), .c(stg2_c1[40]), .co(stg2_co1[40]));
counter_5to3 u_a21_41(.i0(stg1_s1_w[41]), .i1(stg1_c1_w[40]), .i2(stg1_s2_w[33]), .i3(stg1_c2_w[32]), .ci(stg2_co1[40]), .s(stg2_s1[41]), .c(stg2_c1[41]), .co(stg2_co1[41]));
counter_5to3 u_a21_42(.i0(stg1_s1_w[42]), .i1(stg1_c1_w[41]), .i2(stg1_s2_w[34]), .i3(stg1_c2_w[33]), .ci(stg2_co1[41]), .s(stg2_s1[42]), .c(stg2_c1[42]), .co(stg2_co1[42]));
counter_5to3 u_a21_43(.i0(stg1_s1_w[43]), .i1(stg1_c1_w[42]), .i2(stg1_s2_w[35]), .i3(stg1_c2_w[34]), .ci(stg2_co1[42]), .s(stg2_s1[43]), .c(stg2_c1[43]), .co(stg2_co1[43]));
counter_5to3 u_a21_44(.i0(stg1_s1_w[44]), .i1(stg1_c1_w[43]), .i2(stg1_s2_w[36]), .i3(stg1_c2_w[35]), .ci(stg2_co1[43]), .s(stg2_s1[44]), .c(stg2_c1[44]), .co(stg2_co1[44]));
counter_5to3 u_a21_45(.i0(stg1_s1_w[45]), .i1(stg1_c1_w[44]), .i2(stg1_s2_w[37]), .i3(stg1_c2_w[36]), .ci(stg2_co1[44]), .s(stg2_s1[45]), .c(stg2_c1[45]), .co(stg2_co1[45]));
counter_5to3 u_a21_46(.i0(stg1_s1_w[46]), .i1(stg1_c1_w[45]), .i2(stg1_s2_w[38]), .i3(stg1_c2_w[37]), .ci(stg2_co1[45]), .s(stg2_s1[46]), .c(stg2_c1[46]), .co(stg2_co1[46]));
counter_5to3 u_a21_47(.i0(stg1_s1_w[47]), .i1(stg1_c1_w[46]), .i2(stg1_s2_w[39]), .i3(stg1_c2_w[38]), .ci(stg2_co1[46]), .s(stg2_s1[47]), .c(stg2_c1[47]), .co(stg2_co1[47]));
counter_5to3 u_a21_48(.i0(stg1_s1_w[48]), .i1(stg1_c1_w[47]), .i2(stg1_s2_w[40]), .i3(stg1_c2_w[39]), .ci(stg2_co1[47]), .s(stg2_s1[48]), .c(stg2_c1[48]), .co(stg2_co1[48]));
counter_5to3 u_a21_49(.i0(stg1_s1_w[49]), .i1(stg1_c1_w[48]), .i2(stg1_s2_w[41]), .i3(stg1_c2_w[40]), .ci(stg2_co1[48]), .s(stg2_s1[49]), .c(stg2_c1[49]), .co(stg2_co1[49]));
counter_5to3 u_a21_50(.i0(stg1_s1_w[50]), .i1(stg1_c1_w[49]), .i2(stg1_s2_w[42]), .i3(stg1_c2_w[41]), .ci(stg2_co1[49]), .s(stg2_s1[50]), .c(stg2_c1[50]), .co(stg2_co1[50]));
counter_5to3 u_a21_51(.i0(stg1_s1_w[51]), .i1(stg1_c1_w[50]), .i2(stg1_s2_w[43]), .i3(stg1_c2_w[42]), .ci(stg2_co1[50]), .s(stg2_s1[51]), .c(stg2_c1[51]), .co(stg2_co1[51]));
counter_5to3 u_a21_52(.i0(stg1_s1_w[52]), .i1(stg1_c1_w[51]), .i2(stg1_s2_w[44]), .i3(stg1_c2_w[43]), .ci(stg2_co1[51]), .s(stg2_s1[52]), .c(stg2_c1[52]), .co(stg2_co1[52]));
counter_5to3 u_a21_53(.i0(stg1_s1_w[53]), .i1(stg1_c1_w[52]), .i2(stg1_s2_w[45]), .i3(stg1_c2_w[44]), .ci(stg2_co1[52]), .s(stg2_s1[53]), .c(stg2_c1[53]), .co(stg2_co1[53]));
counter_5to3 u_a21_54(.i0(stg1_s1_w[54]), .i1(stg1_c1_w[53]), .i2(stg1_s2_w[46]), .i3(stg1_c2_w[45]), .ci(stg2_co1[53]), .s(stg2_s1[54]), .c(stg2_c1[54]), .co(stg2_co1[54]));
counter_5to3 u_a21_55(.i0(stg1_s1_w[55]), .i1(stg1_c1_w[54]), .i2(stg1_s2_w[47]), .i3(stg1_c2_w[46]), .ci(stg2_co1[54]), .s(stg2_s1[55]), .c(stg2_c1[55]), .co(stg2_co1[55]));
counter_5to3 u_a21_56(.i0(stg1_s1_w[56]), .i1(stg1_c1_w[55]), .i2(stg1_s2_w[48]), .i3(stg1_c2_w[47]), .ci(stg2_co1[55]), .s(stg2_s1[56]), .c(stg2_c1[56]), .co(stg2_co1[56]));
counter_5to3 u_a21_57(.i0(stg1_s1_w[57]), .i1(stg1_c1_w[56]), .i2(stg1_s2_w[49]), .i3(stg1_c2_w[48]), .ci(stg2_co1[56]), .s(stg2_s1[57]), .c(stg2_c1[57]), .co(stg2_co1[57]));
counter_5to3 u_a21_58(.i0(stg1_s1_w[58]), .i1(stg1_c1_w[57]), .i2(stg1_s2_w[50]), .i3(stg1_c2_w[49]), .ci(stg2_co1[57]), .s(stg2_s1[58]), .c(stg2_c1[58]), .co(stg2_co1[58]));
counter_5to3 u_a21_59(.i0(stg1_s1_w[59]), .i1(stg1_c1_w[58]), .i2(stg1_s2_w[51]), .i3(stg1_c2_w[50]), .ci(stg2_co1[58]), .s(stg2_s1[59]), .c(stg2_c1[59]), .co(stg2_co1[59]));
counter_5to3 u_a21_60(.i0(stg1_s1_w[60]), .i1(stg1_c1_w[59]), .i2(stg1_s2_w[52]), .i3(stg1_c2_w[51]), .ci(stg2_co1[59]), .s(stg2_s1[60]), .c(stg2_c1[60]), .co(stg2_co1[60]));
counter_5to3 u_a21_61(.i0(stg1_s1_w[61]), .i1(stg1_c1_w[60]), .i2(stg1_s2_w[53]), .i3(stg1_c2_w[52]), .ci(stg2_co1[60]), .s(stg2_s1[61]), .c(stg2_c1[61]), .co(stg2_co1[61]));
counter_5to3 u_a21_62(.i0(stg1_s1_w[62]), .i1(stg1_c1_w[61]), .i2(stg1_s2_w[54]), .i3(stg1_c2_w[53]), .ci(stg2_co1[61]), .s(stg2_s1[62]), .c(stg2_c1[62]), .co(stg2_co1[62]));
counter_5to3 u_a21_63(.i0(stg1_s1_w[63]), .i1(stg1_c1_w[62]), .i2(stg1_s2_w[55]), .i3(stg1_c2_w[54]), .ci(stg2_co1[62]), .s(stg2_s1[63]), .c(stg2_c1[63]), .co(stg2_co1[63]));
counter_5to3 u_a21_64(.i0(stg1_s1_w[64]), .i1(stg1_c1_w[63]), .i2(stg1_s2_w[56]), .i3(stg1_c2_w[55]), .ci(stg2_co1[63]), .s(stg2_s1[64]), .c(stg2_c1[64]), .co(stg2_co1[64]));
counter_5to3 u_a21_65(.i0(stg1_s1_w[65]), .i1(stg1_c1_w[64]), .i2(stg1_s2_w[57]), .i3(stg1_c2_w[56]), .ci(stg2_co1[64]), .s(stg2_s1[65]), .c(stg2_c1[65]), .co(stg2_co1[65]));
counter_5to3 u_a21_66(.i0(stg1_s1_w[66]), .i1(stg1_c1_w[65]), .i2(stg1_s2_w[58]), .i3(stg1_c2_w[57]), .ci(stg2_co1[65]), .s(stg2_s1[66]), .c(stg2_c1[66]), .co(stg2_co1[66]));
counter_5to3 u_a21_67(.i0(stg1_s1_w[67]), .i1(stg1_c1_w[66]), .i2(stg1_s2_w[59]), .i3(stg1_c2_w[58]), .ci(stg2_co1[66]), .s(stg2_s1[67]), .c(stg2_c1[67]), .co(stg2_co1[67]));
counter_5to3 u_a21_68(.i0(stg1_s1_w[68]), .i1(stg1_c1_w[67]), .i2(stg1_s2_w[60]), .i3(stg1_c2_w[59]), .ci(stg2_co1[67]), .s(stg2_s1[68]), .c(stg2_c1[68]), .co(stg2_co1[68]));
counter_5to3 u_a21_69(.i0(stg1_s1_w[69]), .i1(stg1_c1_w[68]), .i2(stg1_s2_w[61]), .i3(stg1_c2_w[60]), .ci(stg2_co1[68]), .s(stg2_s1[69]), .c(stg2_c1[69]), .co(stg2_co1[69]));
counter_5to3 u_a21_70(.i0(stg1_s1_w[70]), .i1(stg1_c1_w[69]), .i2(stg1_s2_w[62]), .i3(stg1_c2_w[61]), .ci(stg2_co1[69]), .s(stg2_s1[70]), .c(stg2_c1[70]), .co(stg2_co1[70]));
counter_5to3 u_a21_71(.i0(stg1_s1_w[71]), .i1(stg1_c1_w[70]), .i2(stg1_s2_w[63]), .i3(stg1_c2_w[62]), .ci(stg2_co1[70]), .s(stg2_s1[71]), .c(stg2_c1[71]), .co(stg2_co1[71]));
counter_5to3 u_a21_72(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[71]), .i2(stg1_s2_w[64]), .i3(stg1_c2_w[63]), .ci(stg2_co1[71]), .s(stg2_s1[72]), .c(stg2_c1[72]), .co(stg2_co1[72]));
counter_5to3 u_a21_73(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[65]), .i3(stg1_c2_w[64]), .ci(stg2_co1[72]), .s(stg2_s1[73]), .c(stg2_c1[73]), .co(stg2_co1[73]));
counter_5to3 u_a21_74(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[66]), .i3(stg1_c2_w[65]), .ci(stg2_co1[73]), .s(stg2_s1[74]), .c(stg2_c1[74]), .co(stg2_co1[74]));
counter_5to3 u_a21_75(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[67]), .i3(stg1_c2_w[66]), .ci(stg2_co1[74]), .s(stg2_s1[75]), .c(stg2_c1[75]), .co(stg2_co1[75]));
counter_5to3 u_a21_76(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[68]), .i3(stg1_c2_w[67]), .ci(stg2_co1[75]), .s(stg2_s1[76]), .c(stg2_c1[76]), .co(stg2_co1[76]));
counter_5to3 u_a21_77(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[69]), .i3(stg1_c2_w[68]), .ci(stg2_co1[76]), .s(stg2_s1[77]), .c(stg2_c1[77]), .co(stg2_co1[77]));
counter_5to3 u_a21_78(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[70]), .i3(stg1_c2_w[69]), .ci(stg2_co1[77]), .s(stg2_s1[78]), .c(stg2_c1[78]), .co(stg2_co1[78]));
counter_5to3 u_a21_79(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[71]), .i3(stg1_c2_w[70]), .ci(stg2_co1[78]), .s(stg2_s1[79]), .c(stg2_c1[79]), .co(stg2_co1[79]));
counter_5to3 u_a21_80(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[72]), .i3(stg1_c2_w[71]), .ci(stg2_co1[79]), .s(stg2_s1[80]), .c(stg2_c1[80]), .co(stg2_co1[80]));
counter_5to3 u_a21_81(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[72]), .i3(stg1_c2_w[72]), .ci(stg2_co1[80]), .s(stg2_s1[81]), .c(stg2_c1[81]), .co(stg2_co1[81]));
counter_5to3 u_a21_82(.i0(stg1_s1_w[72]), .i1(stg1_c1_w[72]), .i2(stg1_s2_w[72]), .i3(stg1_c2_w[72]), .ci(stg2_co1[81]), .s(stg2_s1[82]), .c(stg2_c1[82]), .co(stg2_co1[82]));

// =========================== second stage 2nd group ============================================================================================================
counter_5to3 u_a22_0 (.i0(stg1_s3_w[0 ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0         ), .ci(1'b0        ), .s(stg2_s2[0 ]), .c(stg2_c2[0 ]), .co(stg2_co2[0 ]));
counter_5to3 u_a22_1 (.i0(stg1_s3_w[1 ]), .i1(stg1_c3_w[0 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[0 ]), .s(stg2_s2[1 ]), .c(stg2_c2[1 ]), .co(stg2_co2[1 ]));
counter_5to3 u_a22_2 (.i0(stg1_s3_w[2 ]), .i1(stg1_c3_w[1 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[1 ]), .s(stg2_s2[2 ]), .c(stg2_c2[2 ]), .co(stg2_co2[2 ]));
counter_5to3 u_a22_3 (.i0(stg1_s3_w[3 ]), .i1(stg1_c3_w[2 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[2 ]), .s(stg2_s2[3 ]), .c(stg2_c2[3 ]), .co(stg2_co2[3 ]));
counter_5to3 u_a22_4 (.i0(stg1_s3_w[4 ]), .i1(stg1_c3_w[3 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[3 ]), .s(stg2_s2[4 ]), .c(stg2_c2[4 ]), .co(stg2_co2[4 ]));
counter_5to3 u_a22_5 (.i0(stg1_s3_w[5 ]), .i1(stg1_c3_w[4 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[4 ]), .s(stg2_s2[5 ]), .c(stg2_c2[5 ]), .co(stg2_co2[5 ]));
counter_5to3 u_a22_6 (.i0(stg1_s3_w[6 ]), .i1(stg1_c3_w[5 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[5 ]), .s(stg2_s2[6 ]), .c(stg2_c2[6 ]), .co(stg2_co2[6 ]));
counter_5to3 u_a22_7 (.i0(stg1_s3_w[7 ]), .i1(stg1_c3_w[6 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co2[6 ]), .s(stg2_s2[7 ]), .c(stg2_c2[7 ]), .co(stg2_co2[7 ]));
counter_5to3 u_a22_8 (.i0(stg1_s3_w[8 ]), .i1(stg1_c3_w[7 ]), .i2(stg1_s4_w[0 ]), .i3(1'b0         ), .ci(stg2_co2[7 ]), .s(stg2_s2[8 ]), .c(stg2_c2[8 ]), .co(stg2_co2[8 ]));
counter_5to3 u_a22_9 (.i0(stg1_s3_w[9 ]), .i1(stg1_c3_w[8 ]), .i2(stg1_s4_w[1 ]), .i3(stg1_c4_w[0 ]), .ci(stg2_co2[8 ]), .s(stg2_s2[9 ]), .c(stg2_c2[9 ]), .co(stg2_co2[9 ]));
counter_5to3 u_a22_10(.i0(stg1_s3_w[10]), .i1(stg1_c3_w[9 ]), .i2(stg1_s4_w[2 ]), .i3(stg1_c4_w[1 ]), .ci(stg2_co2[9 ]), .s(stg2_s2[10]), .c(stg2_c2[10]), .co(stg2_co2[10]));
counter_5to3 u_a22_11(.i0(stg1_s3_w[11]), .i1(stg1_c3_w[10]), .i2(stg1_s4_w[3 ]), .i3(stg1_c4_w[2 ]), .ci(stg2_co2[10]), .s(stg2_s2[11]), .c(stg2_c2[11]), .co(stg2_co2[11]));
counter_5to3 u_a22_12(.i0(stg1_s3_w[12]), .i1(stg1_c3_w[11]), .i2(stg1_s4_w[4 ]), .i3(stg1_c4_w[3 ]), .ci(stg2_co2[11]), .s(stg2_s2[12]), .c(stg2_c2[12]), .co(stg2_co2[12]));
counter_5to3 u_a22_13(.i0(stg1_s3_w[13]), .i1(stg1_c3_w[12]), .i2(stg1_s4_w[5 ]), .i3(stg1_c4_w[4 ]), .ci(stg2_co2[12]), .s(stg2_s2[13]), .c(stg2_c2[13]), .co(stg2_co2[13]));
counter_5to3 u_a22_14(.i0(stg1_s3_w[14]), .i1(stg1_c3_w[13]), .i2(stg1_s4_w[6 ]), .i3(stg1_c4_w[5 ]), .ci(stg2_co2[13]), .s(stg2_s2[14]), .c(stg2_c2[14]), .co(stg2_co2[14]));
counter_5to3 u_a22_15(.i0(stg1_s3_w[15]), .i1(stg1_c3_w[14]), .i2(stg1_s4_w[7 ]), .i3(stg1_c4_w[6 ]), .ci(stg2_co2[14]), .s(stg2_s2[15]), .c(stg2_c2[15]), .co(stg2_co2[15]));
counter_5to3 u_a22_16(.i0(stg1_s3_w[16]), .i1(stg1_c3_w[15]), .i2(stg1_s4_w[8 ]), .i3(stg1_c4_w[7 ]), .ci(stg2_co2[15]), .s(stg2_s2[16]), .c(stg2_c2[16]), .co(stg2_co2[16]));
counter_5to3 u_a22_17(.i0(stg1_s3_w[17]), .i1(stg1_c3_w[16]), .i2(stg1_s4_w[9 ]), .i3(stg1_c4_w[8 ]), .ci(stg2_co2[16]), .s(stg2_s2[17]), .c(stg2_c2[17]), .co(stg2_co2[17]));
counter_5to3 u_a22_18(.i0(stg1_s3_w[18]), .i1(stg1_c3_w[17]), .i2(stg1_s4_w[10]), .i3(stg1_c4_w[9 ]), .ci(stg2_co2[17]), .s(stg2_s2[18]), .c(stg2_c2[18]), .co(stg2_co2[18]));
counter_5to3 u_a22_19(.i0(stg1_s3_w[19]), .i1(stg1_c3_w[18]), .i2(stg1_s4_w[11]), .i3(stg1_c4_w[10]), .ci(stg2_co2[18]), .s(stg2_s2[19]), .c(stg2_c2[19]), .co(stg2_co2[19]));
counter_5to3 u_a22_20(.i0(stg1_s3_w[20]), .i1(stg1_c3_w[19]), .i2(stg1_s4_w[12]), .i3(stg1_c4_w[11]), .ci(stg2_co2[19]), .s(stg2_s2[20]), .c(stg2_c2[20]), .co(stg2_co2[20]));
counter_5to3 u_a22_21(.i0(stg1_s3_w[21]), .i1(stg1_c3_w[20]), .i2(stg1_s4_w[13]), .i3(stg1_c4_w[12]), .ci(stg2_co2[20]), .s(stg2_s2[21]), .c(stg2_c2[21]), .co(stg2_co2[21]));
counter_5to3 u_a22_22(.i0(stg1_s3_w[22]), .i1(stg1_c3_w[21]), .i2(stg1_s4_w[14]), .i3(stg1_c4_w[13]), .ci(stg2_co2[21]), .s(stg2_s2[22]), .c(stg2_c2[22]), .co(stg2_co2[22]));
counter_5to3 u_a22_23(.i0(stg1_s3_w[23]), .i1(stg1_c3_w[22]), .i2(stg1_s4_w[15]), .i3(stg1_c4_w[14]), .ci(stg2_co2[22]), .s(stg2_s2[23]), .c(stg2_c2[23]), .co(stg2_co2[23]));
counter_5to3 u_a22_24(.i0(stg1_s3_w[24]), .i1(stg1_c3_w[23]), .i2(stg1_s4_w[16]), .i3(stg1_c4_w[15]), .ci(stg2_co2[23]), .s(stg2_s2[24]), .c(stg2_c2[24]), .co(stg2_co2[24]));
counter_5to3 u_a22_25(.i0(stg1_s3_w[25]), .i1(stg1_c3_w[24]), .i2(stg1_s4_w[17]), .i3(stg1_c4_w[16]), .ci(stg2_co2[24]), .s(stg2_s2[25]), .c(stg2_c2[25]), .co(stg2_co2[25]));
counter_5to3 u_a22_26(.i0(stg1_s3_w[26]), .i1(stg1_c3_w[25]), .i2(stg1_s4_w[18]), .i3(stg1_c4_w[17]), .ci(stg2_co2[25]), .s(stg2_s2[26]), .c(stg2_c2[26]), .co(stg2_co2[26]));
counter_5to3 u_a22_27(.i0(stg1_s3_w[27]), .i1(stg1_c3_w[26]), .i2(stg1_s4_w[19]), .i3(stg1_c4_w[18]), .ci(stg2_co2[26]), .s(stg2_s2[27]), .c(stg2_c2[27]), .co(stg2_co2[27]));
counter_5to3 u_a22_28(.i0(stg1_s3_w[28]), .i1(stg1_c3_w[27]), .i2(stg1_s4_w[20]), .i3(stg1_c4_w[19]), .ci(stg2_co2[27]), .s(stg2_s2[28]), .c(stg2_c2[28]), .co(stg2_co2[28]));
counter_5to3 u_a22_29(.i0(stg1_s3_w[29]), .i1(stg1_c3_w[28]), .i2(stg1_s4_w[21]), .i3(stg1_c4_w[20]), .ci(stg2_co2[28]), .s(stg2_s2[29]), .c(stg2_c2[29]), .co(stg2_co2[29]));
counter_5to3 u_a22_30(.i0(stg1_s3_w[30]), .i1(stg1_c3_w[29]), .i2(stg1_s4_w[22]), .i3(stg1_c4_w[21]), .ci(stg2_co2[29]), .s(stg2_s2[30]), .c(stg2_c2[30]), .co(stg2_co2[30]));
counter_5to3 u_a22_31(.i0(stg1_s3_w[31]), .i1(stg1_c3_w[30]), .i2(stg1_s4_w[23]), .i3(stg1_c4_w[22]), .ci(stg2_co2[30]), .s(stg2_s2[31]), .c(stg2_c2[31]), .co(stg2_co2[31]));
counter_5to3 u_a22_32(.i0(stg1_s3_w[32]), .i1(stg1_c3_w[31]), .i2(stg1_s4_w[24]), .i3(stg1_c4_w[23]), .ci(stg2_co2[31]), .s(stg2_s2[32]), .c(stg2_c2[32]), .co(stg2_co2[32]));
counter_5to3 u_a22_33(.i0(stg1_s3_w[33]), .i1(stg1_c3_w[32]), .i2(stg1_s4_w[25]), .i3(stg1_c4_w[24]), .ci(stg2_co2[32]), .s(stg2_s2[33]), .c(stg2_c2[33]), .co(stg2_co2[33]));
counter_5to3 u_a22_34(.i0(stg1_s3_w[34]), .i1(stg1_c3_w[33]), .i2(stg1_s4_w[26]), .i3(stg1_c4_w[25]), .ci(stg2_co2[33]), .s(stg2_s2[34]), .c(stg2_c2[34]), .co(stg2_co2[34]));
counter_5to3 u_a22_35(.i0(stg1_s3_w[35]), .i1(stg1_c3_w[34]), .i2(stg1_s4_w[27]), .i3(stg1_c4_w[26]), .ci(stg2_co2[34]), .s(stg2_s2[35]), .c(stg2_c2[35]), .co(stg2_co2[35]));
counter_5to3 u_a22_36(.i0(stg1_s3_w[36]), .i1(stg1_c3_w[35]), .i2(stg1_s4_w[28]), .i3(stg1_c4_w[27]), .ci(stg2_co2[35]), .s(stg2_s2[36]), .c(stg2_c2[36]), .co(stg2_co2[36]));
counter_5to3 u_a22_37(.i0(stg1_s3_w[37]), .i1(stg1_c3_w[36]), .i2(stg1_s4_w[29]), .i3(stg1_c4_w[28]), .ci(stg2_co2[36]), .s(stg2_s2[37]), .c(stg2_c2[37]), .co(stg2_co2[37]));
counter_5to3 u_a22_38(.i0(stg1_s3_w[38]), .i1(stg1_c3_w[37]), .i2(stg1_s4_w[30]), .i3(stg1_c4_w[29]), .ci(stg2_co2[37]), .s(stg2_s2[38]), .c(stg2_c2[38]), .co(stg2_co2[38]));
counter_5to3 u_a22_39(.i0(stg1_s3_w[39]), .i1(stg1_c3_w[38]), .i2(stg1_s4_w[31]), .i3(stg1_c4_w[30]), .ci(stg2_co2[38]), .s(stg2_s2[39]), .c(stg2_c2[39]), .co(stg2_co2[39]));
counter_5to3 u_a22_40(.i0(stg1_s3_w[40]), .i1(stg1_c3_w[39]), .i2(stg1_s4_w[32]), .i3(stg1_c4_w[31]), .ci(stg2_co2[39]), .s(stg2_s2[40]), .c(stg2_c2[40]), .co(stg2_co2[40]));
counter_5to3 u_a22_41(.i0(stg1_s3_w[41]), .i1(stg1_c3_w[40]), .i2(stg1_s4_w[33]), .i3(stg1_c4_w[32]), .ci(stg2_co2[40]), .s(stg2_s2[41]), .c(stg2_c2[41]), .co(stg2_co2[41]));
counter_5to3 u_a22_42(.i0(stg1_s3_w[42]), .i1(stg1_c3_w[41]), .i2(stg1_s4_w[34]), .i3(stg1_c4_w[33]), .ci(stg2_co2[41]), .s(stg2_s2[42]), .c(stg2_c2[42]), .co(stg2_co2[42]));
counter_5to3 u_a22_43(.i0(stg1_s3_w[43]), .i1(stg1_c3_w[42]), .i2(stg1_s4_w[35]), .i3(stg1_c4_w[34]), .ci(stg2_co2[42]), .s(stg2_s2[43]), .c(stg2_c2[43]), .co(stg2_co2[43]));
counter_5to3 u_a22_44(.i0(stg1_s3_w[44]), .i1(stg1_c3_w[43]), .i2(stg1_s4_w[36]), .i3(stg1_c4_w[35]), .ci(stg2_co2[43]), .s(stg2_s2[44]), .c(stg2_c2[44]), .co(stg2_co2[44]));
counter_5to3 u_a22_45(.i0(stg1_s3_w[45]), .i1(stg1_c3_w[44]), .i2(stg1_s4_w[37]), .i3(stg1_c4_w[36]), .ci(stg2_co2[44]), .s(stg2_s2[45]), .c(stg2_c2[45]), .co(stg2_co2[45]));
counter_5to3 u_a22_46(.i0(stg1_s3_w[46]), .i1(stg1_c3_w[45]), .i2(stg1_s4_w[38]), .i3(stg1_c4_w[37]), .ci(stg2_co2[45]), .s(stg2_s2[46]), .c(stg2_c2[46]), .co(stg2_co2[46]));
counter_5to3 u_a22_47(.i0(stg1_s3_w[47]), .i1(stg1_c3_w[46]), .i2(stg1_s4_w[39]), .i3(stg1_c4_w[38]), .ci(stg2_co2[46]), .s(stg2_s2[47]), .c(stg2_c2[47]), .co(stg2_co2[47]));
counter_5to3 u_a22_48(.i0(stg1_s3_w[48]), .i1(stg1_c3_w[47]), .i2(stg1_s4_w[40]), .i3(stg1_c4_w[39]), .ci(stg2_co2[47]), .s(stg2_s2[48]), .c(stg2_c2[48]), .co(stg2_co2[48]));
counter_5to3 u_a22_49(.i0(stg1_s3_w[49]), .i1(stg1_c3_w[48]), .i2(stg1_s4_w[41]), .i3(stg1_c4_w[40]), .ci(stg2_co2[48]), .s(stg2_s2[49]), .c(stg2_c2[49]), .co(stg2_co2[49]));
counter_5to3 u_a22_50(.i0(stg1_s3_w[50]), .i1(stg1_c3_w[49]), .i2(stg1_s4_w[42]), .i3(stg1_c4_w[41]), .ci(stg2_co2[49]), .s(stg2_s2[50]), .c(stg2_c2[50]), .co(stg2_co2[50]));
counter_5to3 u_a22_51(.i0(stg1_s3_w[51]), .i1(stg1_c3_w[50]), .i2(stg1_s4_w[43]), .i3(stg1_c4_w[42]), .ci(stg2_co2[50]), .s(stg2_s2[51]), .c(stg2_c2[51]), .co(stg2_co2[51]));
counter_5to3 u_a22_52(.i0(stg1_s3_w[52]), .i1(stg1_c3_w[51]), .i2(stg1_s4_w[44]), .i3(stg1_c4_w[43]), .ci(stg2_co2[51]), .s(stg2_s2[52]), .c(stg2_c2[52]), .co(stg2_co2[52]));
counter_5to3 u_a22_53(.i0(stg1_s3_w[53]), .i1(stg1_c3_w[52]), .i2(stg1_s4_w[45]), .i3(stg1_c4_w[44]), .ci(stg2_co2[52]), .s(stg2_s2[53]), .c(stg2_c2[53]), .co(stg2_co2[53]));
counter_5to3 u_a22_54(.i0(stg1_s3_w[54]), .i1(stg1_c3_w[53]), .i2(stg1_s4_w[46]), .i3(stg1_c4_w[45]), .ci(stg2_co2[53]), .s(stg2_s2[54]), .c(stg2_c2[54]), .co(stg2_co2[54]));
counter_5to3 u_a22_55(.i0(stg1_s3_w[55]), .i1(stg1_c3_w[54]), .i2(stg1_s4_w[47]), .i3(stg1_c4_w[46]), .ci(stg2_co2[54]), .s(stg2_s2[55]), .c(stg2_c2[55]), .co(stg2_co2[55]));
counter_5to3 u_a22_56(.i0(stg1_s3_w[56]), .i1(stg1_c3_w[55]), .i2(stg1_s4_w[48]), .i3(stg1_c4_w[47]), .ci(stg2_co2[55]), .s(stg2_s2[56]), .c(stg2_c2[56]), .co(stg2_co2[56]));
counter_5to3 u_a22_57(.i0(stg1_s3_w[57]), .i1(stg1_c3_w[56]), .i2(stg1_s4_w[49]), .i3(stg1_c4_w[48]), .ci(stg2_co2[56]), .s(stg2_s2[57]), .c(stg2_c2[57]), .co(stg2_co2[57]));
counter_5to3 u_a22_58(.i0(stg1_s3_w[58]), .i1(stg1_c3_w[57]), .i2(stg1_s4_w[50]), .i3(stg1_c4_w[49]), .ci(stg2_co2[57]), .s(stg2_s2[58]), .c(stg2_c2[58]), .co(stg2_co2[58]));
counter_5to3 u_a22_59(.i0(stg1_s3_w[59]), .i1(stg1_c3_w[58]), .i2(stg1_s4_w[51]), .i3(stg1_c4_w[50]), .ci(stg2_co2[58]), .s(stg2_s2[59]), .c(stg2_c2[59]), .co(stg2_co2[59]));
counter_5to3 u_a22_60(.i0(stg1_s3_w[60]), .i1(stg1_c3_w[59]), .i2(stg1_s4_w[52]), .i3(stg1_c4_w[51]), .ci(stg2_co2[59]), .s(stg2_s2[60]), .c(stg2_c2[60]), .co(stg2_co2[60]));
counter_5to3 u_a22_61(.i0(stg1_s3_w[61]), .i1(stg1_c3_w[60]), .i2(stg1_s4_w[53]), .i3(stg1_c4_w[52]), .ci(stg2_co2[60]), .s(stg2_s2[61]), .c(stg2_c2[61]), .co(stg2_co2[61]));
counter_5to3 u_a22_62(.i0(stg1_s3_w[62]), .i1(stg1_c3_w[61]), .i2(stg1_s4_w[54]), .i3(stg1_c4_w[53]), .ci(stg2_co2[61]), .s(stg2_s2[62]), .c(stg2_c2[62]), .co(stg2_co2[62]));
counter_5to3 u_a22_63(.i0(stg1_s3_w[63]), .i1(stg1_c3_w[62]), .i2(stg1_s4_w[55]), .i3(stg1_c4_w[54]), .ci(stg2_co2[62]), .s(stg2_s2[63]), .c(stg2_c2[63]), .co(stg2_co2[63]));
counter_5to3 u_a22_64(.i0(stg1_s3_w[64]), .i1(stg1_c3_w[63]), .i2(stg1_s4_w[56]), .i3(stg1_c4_w[55]), .ci(stg2_co2[63]), .s(stg2_s2[64]), .c(stg2_c2[64]), .co(stg2_co2[64]));
counter_5to3 u_a22_65(.i0(stg1_s3_w[65]), .i1(stg1_c3_w[64]), .i2(stg1_s4_w[57]), .i3(stg1_c4_w[56]), .ci(stg2_co2[64]), .s(stg2_s2[65]), .c(stg2_c2[65]), .co(stg2_co2[65]));
counter_5to3 u_a22_66(.i0(stg1_s3_w[66]), .i1(stg1_c3_w[65]), .i2(stg1_s4_w[58]), .i3(stg1_c4_w[57]), .ci(stg2_co2[65]), .s(stg2_s2[66]), .c(stg2_c2[66]), .co(stg2_co2[66]));
counter_5to3 u_a22_67(.i0(stg1_s3_w[67]), .i1(stg1_c3_w[66]), .i2(stg1_s4_w[59]), .i3(stg1_c4_w[58]), .ci(stg2_co2[66]), .s(stg2_s2[67]), .c(stg2_c2[67]), .co(stg2_co2[67]));
counter_5to3 u_a22_68(.i0(stg1_s3_w[68]), .i1(stg1_c3_w[67]), .i2(stg1_s4_w[60]), .i3(stg1_c4_w[59]), .ci(stg2_co2[67]), .s(stg2_s2[68]), .c(stg2_c2[68]), .co(stg2_co2[68]));
counter_5to3 u_a22_69(.i0(stg1_s3_w[69]), .i1(stg1_c3_w[68]), .i2(stg1_s4_w[61]), .i3(stg1_c4_w[60]), .ci(stg2_co2[68]), .s(stg2_s2[69]), .c(stg2_c2[69]), .co(stg2_co2[69]));
counter_5to3 u_a22_70(.i0(stg1_s3_w[70]), .i1(stg1_c3_w[69]), .i2(stg1_s4_w[62]), .i3(stg1_c4_w[61]), .ci(stg2_co2[69]), .s(stg2_s2[70]), .c(stg2_c2[70]), .co(stg2_co2[70]));
counter_5to3 u_a22_71(.i0(stg1_s3_w[71]), .i1(stg1_c3_w[70]), .i2(stg1_s4_w[63]), .i3(stg1_c4_w[62]), .ci(stg2_co2[70]), .s(stg2_s2[71]), .c(stg2_c2[71]), .co(stg2_co2[71]));
counter_5to3 u_a22_72(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[71]), .i2(stg1_s4_w[64]), .i3(stg1_c4_w[63]), .ci(stg2_co2[71]), .s(stg2_s2[72]), .c(stg2_c2[72]), .co(stg2_co2[72]));
counter_5to3 u_a22_73(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[65]), .i3(stg1_c4_w[64]), .ci(stg2_co2[72]), .s(stg2_s2[73]), .c(stg2_c2[73]), .co(stg2_co2[73]));
counter_5to3 u_a22_74(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[66]), .i3(stg1_c4_w[65]), .ci(stg2_co2[73]), .s(stg2_s2[74]), .c(stg2_c2[74]), .co(stg2_co2[74]));
counter_5to3 u_a22_75(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[67]), .i3(stg1_c4_w[66]), .ci(stg2_co2[74]), .s(stg2_s2[75]), .c(stg2_c2[75]), .co(stg2_co2[75]));
counter_5to3 u_a22_76(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[68]), .i3(stg1_c4_w[67]), .ci(stg2_co2[75]), .s(stg2_s2[76]), .c(stg2_c2[76]), .co(stg2_co2[76]));
counter_5to3 u_a22_77(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[69]), .i3(stg1_c4_w[68]), .ci(stg2_co2[76]), .s(stg2_s2[77]), .c(stg2_c2[77]), .co(stg2_co2[77]));
counter_5to3 u_a22_78(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[70]), .i3(stg1_c4_w[69]), .ci(stg2_co2[77]), .s(stg2_s2[78]), .c(stg2_c2[78]), .co(stg2_co2[78]));
counter_5to3 u_a22_79(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[71]), .i3(stg1_c4_w[70]), .ci(stg2_co2[78]), .s(stg2_s2[79]), .c(stg2_c2[79]), .co(stg2_co2[79]));
counter_5to3 u_a22_80(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[72]), .i3(stg1_c4_w[71]), .ci(stg2_co2[79]), .s(stg2_s2[80]), .c(stg2_c2[80]), .co(stg2_co2[80]));
counter_5to3 u_a22_81(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[72]), .i3(stg1_c4_w[72]), .ci(stg2_co2[80]), .s(stg2_s2[81]), .c(stg2_c2[81]), .co(stg2_co2[81]));
counter_5to3 u_a22_82(.i0(stg1_s3_w[72]), .i1(stg1_c3_w[72]), .i2(stg1_s4_w[72]), .i3(stg1_c4_w[72]), .ci(stg2_co2[81]), .s(stg2_s2[82]), .c(stg2_c2[82]), .co(stg2_co2[82]));

// =========================== second stage 3rd group ============================================================================================================
counter_5to3 u_a23_0 (.i0(stg1_s5_w[0 ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0         ), .ci(1'b0        ), .s(stg2_s3[0 ]), .c(stg2_c3[0 ]), .co(stg2_co3[0 ]));
counter_5to3 u_a23_1 (.i0(stg1_s5_w[1 ]), .i1(stg1_c5_w[0 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[0 ]), .s(stg2_s3[1 ]), .c(stg2_c3[1 ]), .co(stg2_co3[1 ]));
counter_5to3 u_a23_2 (.i0(stg1_s5_w[2 ]), .i1(stg1_c5_w[1 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[1 ]), .s(stg2_s3[2 ]), .c(stg2_c3[2 ]), .co(stg2_co3[2 ]));
counter_5to3 u_a23_3 (.i0(stg1_s5_w[3 ]), .i1(stg1_c5_w[2 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[2 ]), .s(stg2_s3[3 ]), .c(stg2_c3[3 ]), .co(stg2_co3[3 ]));
counter_5to3 u_a23_4 (.i0(stg1_s5_w[4 ]), .i1(stg1_c5_w[3 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[3 ]), .s(stg2_s3[4 ]), .c(stg2_c3[4 ]), .co(stg2_co3[4 ]));
counter_5to3 u_a23_5 (.i0(stg1_s5_w[5 ]), .i1(stg1_c5_w[4 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[4 ]), .s(stg2_s3[5 ]), .c(stg2_c3[5 ]), .co(stg2_co3[5 ]));
counter_5to3 u_a23_6 (.i0(stg1_s5_w[6 ]), .i1(stg1_c5_w[5 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[5 ]), .s(stg2_s3[6 ]), .c(stg2_c3[6 ]), .co(stg2_co3[6 ]));
counter_5to3 u_a23_7 (.i0(stg1_s5_w[7 ]), .i1(stg1_c5_w[6 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co3[6 ]), .s(stg2_s3[7 ]), .c(stg2_c3[7 ]), .co(stg2_co3[7 ]));
counter_5to3 u_a23_8 (.i0(stg1_s5_w[8 ]), .i1(stg1_c5_w[7 ]), .i2(stg1_s6_w[0 ]), .i3(1'b0         ), .ci(stg2_co3[7 ]), .s(stg2_s3[8 ]), .c(stg2_c3[8 ]), .co(stg2_co3[8 ]));
counter_5to3 u_a23_9 (.i0(stg1_s5_w[9 ]), .i1(stg1_c5_w[8 ]), .i2(stg1_s6_w[1 ]), .i3(stg1_c6_w[0 ]), .ci(stg2_co3[8 ]), .s(stg2_s3[9 ]), .c(stg2_c3[9 ]), .co(stg2_co3[9 ]));
counter_5to3 u_a23_10(.i0(stg1_s5_w[10]), .i1(stg1_c5_w[9 ]), .i2(stg1_s6_w[2 ]), .i3(stg1_c6_w[1 ]), .ci(stg2_co3[9 ]), .s(stg2_s3[10]), .c(stg2_c3[10]), .co(stg2_co3[10]));
counter_5to3 u_a23_11(.i0(stg1_s5_w[11]), .i1(stg1_c5_w[10]), .i2(stg1_s6_w[3 ]), .i3(stg1_c6_w[2 ]), .ci(stg2_co3[10]), .s(stg2_s3[11]), .c(stg2_c3[11]), .co(stg2_co3[11]));
counter_5to3 u_a23_12(.i0(stg1_s5_w[12]), .i1(stg1_c5_w[11]), .i2(stg1_s6_w[4 ]), .i3(stg1_c6_w[3 ]), .ci(stg2_co3[11]), .s(stg2_s3[12]), .c(stg2_c3[12]), .co(stg2_co3[12]));
counter_5to3 u_a23_13(.i0(stg1_s5_w[13]), .i1(stg1_c5_w[12]), .i2(stg1_s6_w[5 ]), .i3(stg1_c6_w[4 ]), .ci(stg2_co3[12]), .s(stg2_s3[13]), .c(stg2_c3[13]), .co(stg2_co3[13]));
counter_5to3 u_a23_14(.i0(stg1_s5_w[14]), .i1(stg1_c5_w[13]), .i2(stg1_s6_w[6 ]), .i3(stg1_c6_w[5 ]), .ci(stg2_co3[13]), .s(stg2_s3[14]), .c(stg2_c3[14]), .co(stg2_co3[14]));
counter_5to3 u_a23_15(.i0(stg1_s5_w[15]), .i1(stg1_c5_w[14]), .i2(stg1_s6_w[7 ]), .i3(stg1_c6_w[6 ]), .ci(stg2_co3[14]), .s(stg2_s3[15]), .c(stg2_c3[15]), .co(stg2_co3[15]));
counter_5to3 u_a23_16(.i0(stg1_s5_w[16]), .i1(stg1_c5_w[15]), .i2(stg1_s6_w[8 ]), .i3(stg1_c6_w[7 ]), .ci(stg2_co3[15]), .s(stg2_s3[16]), .c(stg2_c3[16]), .co(stg2_co3[16]));
counter_5to3 u_a23_17(.i0(stg1_s5_w[17]), .i1(stg1_c5_w[16]), .i2(stg1_s6_w[9 ]), .i3(stg1_c6_w[8 ]), .ci(stg2_co3[16]), .s(stg2_s3[17]), .c(stg2_c3[17]), .co(stg2_co3[17]));
counter_5to3 u_a23_18(.i0(stg1_s5_w[18]), .i1(stg1_c5_w[17]), .i2(stg1_s6_w[10]), .i3(stg1_c6_w[9 ]), .ci(stg2_co3[17]), .s(stg2_s3[18]), .c(stg2_c3[18]), .co(stg2_co3[18]));
counter_5to3 u_a23_19(.i0(stg1_s5_w[19]), .i1(stg1_c5_w[18]), .i2(stg1_s6_w[11]), .i3(stg1_c6_w[10]), .ci(stg2_co3[18]), .s(stg2_s3[19]), .c(stg2_c3[19]), .co(stg2_co3[19]));
counter_5to3 u_a23_20(.i0(stg1_s5_w[20]), .i1(stg1_c5_w[19]), .i2(stg1_s6_w[12]), .i3(stg1_c6_w[11]), .ci(stg2_co3[19]), .s(stg2_s3[20]), .c(stg2_c3[20]), .co(stg2_co3[20]));
counter_5to3 u_a23_21(.i0(stg1_s5_w[21]), .i1(stg1_c5_w[20]), .i2(stg1_s6_w[13]), .i3(stg1_c6_w[12]), .ci(stg2_co3[20]), .s(stg2_s3[21]), .c(stg2_c3[21]), .co(stg2_co3[21]));
counter_5to3 u_a23_22(.i0(stg1_s5_w[22]), .i1(stg1_c5_w[21]), .i2(stg1_s6_w[14]), .i3(stg1_c6_w[13]), .ci(stg2_co3[21]), .s(stg2_s3[22]), .c(stg2_c3[22]), .co(stg2_co3[22]));
counter_5to3 u_a23_23(.i0(stg1_s5_w[23]), .i1(stg1_c5_w[22]), .i2(stg1_s6_w[15]), .i3(stg1_c6_w[14]), .ci(stg2_co3[22]), .s(stg2_s3[23]), .c(stg2_c3[23]), .co(stg2_co3[23]));
counter_5to3 u_a23_24(.i0(stg1_s5_w[24]), .i1(stg1_c5_w[23]), .i2(stg1_s6_w[16]), .i3(stg1_c6_w[15]), .ci(stg2_co3[23]), .s(stg2_s3[24]), .c(stg2_c3[24]), .co(stg2_co3[24]));
counter_5to3 u_a23_25(.i0(stg1_s5_w[25]), .i1(stg1_c5_w[24]), .i2(stg1_s6_w[17]), .i3(stg1_c6_w[16]), .ci(stg2_co3[24]), .s(stg2_s3[25]), .c(stg2_c3[25]), .co(stg2_co3[25]));
counter_5to3 u_a23_26(.i0(stg1_s5_w[26]), .i1(stg1_c5_w[25]), .i2(stg1_s6_w[18]), .i3(stg1_c6_w[17]), .ci(stg2_co3[25]), .s(stg2_s3[26]), .c(stg2_c3[26]), .co(stg2_co3[26]));
counter_5to3 u_a23_27(.i0(stg1_s5_w[27]), .i1(stg1_c5_w[26]), .i2(stg1_s6_w[19]), .i3(stg1_c6_w[18]), .ci(stg2_co3[26]), .s(stg2_s3[27]), .c(stg2_c3[27]), .co(stg2_co3[27]));
counter_5to3 u_a23_28(.i0(stg1_s5_w[28]), .i1(stg1_c5_w[27]), .i2(stg1_s6_w[20]), .i3(stg1_c6_w[19]), .ci(stg2_co3[27]), .s(stg2_s3[28]), .c(stg2_c3[28]), .co(stg2_co3[28]));
counter_5to3 u_a23_29(.i0(stg1_s5_w[29]), .i1(stg1_c5_w[28]), .i2(stg1_s6_w[21]), .i3(stg1_c6_w[20]), .ci(stg2_co3[28]), .s(stg2_s3[29]), .c(stg2_c3[29]), .co(stg2_co3[29]));
counter_5to3 u_a23_30(.i0(stg1_s5_w[30]), .i1(stg1_c5_w[29]), .i2(stg1_s6_w[22]), .i3(stg1_c6_w[21]), .ci(stg2_co3[29]), .s(stg2_s3[30]), .c(stg2_c3[30]), .co(stg2_co3[30]));
counter_5to3 u_a23_31(.i0(stg1_s5_w[31]), .i1(stg1_c5_w[30]), .i2(stg1_s6_w[23]), .i3(stg1_c6_w[22]), .ci(stg2_co3[30]), .s(stg2_s3[31]), .c(stg2_c3[31]), .co(stg2_co3[31]));
counter_5to3 u_a23_32(.i0(stg1_s5_w[32]), .i1(stg1_c5_w[31]), .i2(stg1_s6_w[24]), .i3(stg1_c6_w[23]), .ci(stg2_co3[31]), .s(stg2_s3[32]), .c(stg2_c3[32]), .co(stg2_co3[32]));
counter_5to3 u_a23_33(.i0(stg1_s5_w[33]), .i1(stg1_c5_w[32]), .i2(stg1_s6_w[25]), .i3(stg1_c6_w[24]), .ci(stg2_co3[32]), .s(stg2_s3[33]), .c(stg2_c3[33]), .co(stg2_co3[33]));
counter_5to3 u_a23_34(.i0(stg1_s5_w[34]), .i1(stg1_c5_w[33]), .i2(stg1_s6_w[26]), .i3(stg1_c6_w[25]), .ci(stg2_co3[33]), .s(stg2_s3[34]), .c(stg2_c3[34]), .co(stg2_co3[34]));
counter_5to3 u_a23_35(.i0(stg1_s5_w[35]), .i1(stg1_c5_w[34]), .i2(stg1_s6_w[27]), .i3(stg1_c6_w[26]), .ci(stg2_co3[34]), .s(stg2_s3[35]), .c(stg2_c3[35]), .co(stg2_co3[35]));
counter_5to3 u_a23_36(.i0(stg1_s5_w[36]), .i1(stg1_c5_w[35]), .i2(stg1_s6_w[28]), .i3(stg1_c6_w[27]), .ci(stg2_co3[35]), .s(stg2_s3[36]), .c(stg2_c3[36]), .co(stg2_co3[36]));
counter_5to3 u_a23_37(.i0(stg1_s5_w[37]), .i1(stg1_c5_w[36]), .i2(stg1_s6_w[29]), .i3(stg1_c6_w[28]), .ci(stg2_co3[36]), .s(stg2_s3[37]), .c(stg2_c3[37]), .co(stg2_co3[37]));
counter_5to3 u_a23_38(.i0(stg1_s5_w[38]), .i1(stg1_c5_w[37]), .i2(stg1_s6_w[30]), .i3(stg1_c6_w[29]), .ci(stg2_co3[37]), .s(stg2_s3[38]), .c(stg2_c3[38]), .co(stg2_co3[38]));
counter_5to3 u_a23_39(.i0(stg1_s5_w[39]), .i1(stg1_c5_w[38]), .i2(stg1_s6_w[31]), .i3(stg1_c6_w[30]), .ci(stg2_co3[38]), .s(stg2_s3[39]), .c(stg2_c3[39]), .co(stg2_co3[39]));
counter_5to3 u_a23_40(.i0(stg1_s5_w[40]), .i1(stg1_c5_w[39]), .i2(stg1_s6_w[32]), .i3(stg1_c6_w[31]), .ci(stg2_co3[39]), .s(stg2_s3[40]), .c(stg2_c3[40]), .co(stg2_co3[40]));
counter_5to3 u_a23_41(.i0(stg1_s5_w[41]), .i1(stg1_c5_w[40]), .i2(stg1_s6_w[33]), .i3(stg1_c6_w[32]), .ci(stg2_co3[40]), .s(stg2_s3[41]), .c(stg2_c3[41]), .co(stg2_co3[41]));
counter_5to3 u_a23_42(.i0(stg1_s5_w[42]), .i1(stg1_c5_w[41]), .i2(stg1_s6_w[34]), .i3(stg1_c6_w[33]), .ci(stg2_co3[41]), .s(stg2_s3[42]), .c(stg2_c3[42]), .co(stg2_co3[42]));
counter_5to3 u_a23_43(.i0(stg1_s5_w[43]), .i1(stg1_c5_w[42]), .i2(stg1_s6_w[35]), .i3(stg1_c6_w[34]), .ci(stg2_co3[42]), .s(stg2_s3[43]), .c(stg2_c3[43]), .co(stg2_co3[43]));
counter_5to3 u_a23_44(.i0(stg1_s5_w[44]), .i1(stg1_c5_w[43]), .i2(stg1_s6_w[36]), .i3(stg1_c6_w[35]), .ci(stg2_co3[43]), .s(stg2_s3[44]), .c(stg2_c3[44]), .co(stg2_co3[44]));
counter_5to3 u_a23_45(.i0(stg1_s5_w[45]), .i1(stg1_c5_w[44]), .i2(stg1_s6_w[37]), .i3(stg1_c6_w[36]), .ci(stg2_co3[44]), .s(stg2_s3[45]), .c(stg2_c3[45]), .co(stg2_co3[45]));
counter_5to3 u_a23_46(.i0(stg1_s5_w[46]), .i1(stg1_c5_w[45]), .i2(stg1_s6_w[38]), .i3(stg1_c6_w[37]), .ci(stg2_co3[45]), .s(stg2_s3[46]), .c(stg2_c3[46]), .co(stg2_co3[46]));
counter_5to3 u_a23_47(.i0(stg1_s5_w[47]), .i1(stg1_c5_w[46]), .i2(stg1_s6_w[39]), .i3(stg1_c6_w[38]), .ci(stg2_co3[46]), .s(stg2_s3[47]), .c(stg2_c3[47]), .co(stg2_co3[47]));
counter_5to3 u_a23_48(.i0(stg1_s5_w[48]), .i1(stg1_c5_w[47]), .i2(stg1_s6_w[40]), .i3(stg1_c6_w[39]), .ci(stg2_co3[47]), .s(stg2_s3[48]), .c(stg2_c3[48]), .co(stg2_co3[48]));
counter_5to3 u_a23_49(.i0(stg1_s5_w[49]), .i1(stg1_c5_w[48]), .i2(stg1_s6_w[41]), .i3(stg1_c6_w[40]), .ci(stg2_co3[48]), .s(stg2_s3[49]), .c(stg2_c3[49]), .co(stg2_co3[49]));
counter_5to3 u_a23_50(.i0(stg1_s5_w[50]), .i1(stg1_c5_w[49]), .i2(stg1_s6_w[42]), .i3(stg1_c6_w[41]), .ci(stg2_co3[49]), .s(stg2_s3[50]), .c(stg2_c3[50]), .co(stg2_co3[50]));
counter_5to3 u_a23_51(.i0(stg1_s5_w[51]), .i1(stg1_c5_w[50]), .i2(stg1_s6_w[43]), .i3(stg1_c6_w[42]), .ci(stg2_co3[50]), .s(stg2_s3[51]), .c(stg2_c3[51]), .co(stg2_co3[51]));
counter_5to3 u_a23_52(.i0(stg1_s5_w[52]), .i1(stg1_c5_w[51]), .i2(stg1_s6_w[44]), .i3(stg1_c6_w[43]), .ci(stg2_co3[51]), .s(stg2_s3[52]), .c(stg2_c3[52]), .co(stg2_co3[52]));
counter_5to3 u_a23_53(.i0(stg1_s5_w[53]), .i1(stg1_c5_w[52]), .i2(stg1_s6_w[45]), .i3(stg1_c6_w[44]), .ci(stg2_co3[52]), .s(stg2_s3[53]), .c(stg2_c3[53]), .co(stg2_co3[53]));
counter_5to3 u_a23_54(.i0(stg1_s5_w[54]), .i1(stg1_c5_w[53]), .i2(stg1_s6_w[46]), .i3(stg1_c6_w[45]), .ci(stg2_co3[53]), .s(stg2_s3[54]), .c(stg2_c3[54]), .co(stg2_co3[54]));
counter_5to3 u_a23_55(.i0(stg1_s5_w[55]), .i1(stg1_c5_w[54]), .i2(stg1_s6_w[47]), .i3(stg1_c6_w[46]), .ci(stg2_co3[54]), .s(stg2_s3[55]), .c(stg2_c3[55]), .co(stg2_co3[55]));
counter_5to3 u_a23_56(.i0(stg1_s5_w[56]), .i1(stg1_c5_w[55]), .i2(stg1_s6_w[48]), .i3(stg1_c6_w[47]), .ci(stg2_co3[55]), .s(stg2_s3[56]), .c(stg2_c3[56]), .co(stg2_co3[56]));
counter_5to3 u_a23_57(.i0(stg1_s5_w[57]), .i1(stg1_c5_w[56]), .i2(stg1_s6_w[49]), .i3(stg1_c6_w[48]), .ci(stg2_co3[56]), .s(stg2_s3[57]), .c(stg2_c3[57]), .co(stg2_co3[57]));
counter_5to3 u_a23_58(.i0(stg1_s5_w[58]), .i1(stg1_c5_w[57]), .i2(stg1_s6_w[50]), .i3(stg1_c6_w[49]), .ci(stg2_co3[57]), .s(stg2_s3[58]), .c(stg2_c3[58]), .co(stg2_co3[58]));
counter_5to3 u_a23_59(.i0(stg1_s5_w[59]), .i1(stg1_c5_w[58]), .i2(stg1_s6_w[51]), .i3(stg1_c6_w[50]), .ci(stg2_co3[58]), .s(stg2_s3[59]), .c(stg2_c3[59]), .co(stg2_co3[59]));
counter_5to3 u_a23_60(.i0(stg1_s5_w[60]), .i1(stg1_c5_w[59]), .i2(stg1_s6_w[52]), .i3(stg1_c6_w[51]), .ci(stg2_co3[59]), .s(stg2_s3[60]), .c(stg2_c3[60]), .co(stg2_co3[60]));
counter_5to3 u_a23_61(.i0(stg1_s5_w[61]), .i1(stg1_c5_w[60]), .i2(stg1_s6_w[53]), .i3(stg1_c6_w[52]), .ci(stg2_co3[60]), .s(stg2_s3[61]), .c(stg2_c3[61]), .co(stg2_co3[61]));
counter_5to3 u_a23_62(.i0(stg1_s5_w[62]), .i1(stg1_c5_w[61]), .i2(stg1_s6_w[54]), .i3(stg1_c6_w[53]), .ci(stg2_co3[61]), .s(stg2_s3[62]), .c(stg2_c3[62]), .co(stg2_co3[62]));
counter_5to3 u_a23_63(.i0(stg1_s5_w[63]), .i1(stg1_c5_w[62]), .i2(stg1_s6_w[55]), .i3(stg1_c6_w[54]), .ci(stg2_co3[62]), .s(stg2_s3[63]), .c(stg2_c3[63]), .co(stg2_co3[63]));
counter_5to3 u_a23_64(.i0(stg1_s5_w[64]), .i1(stg1_c5_w[63]), .i2(stg1_s6_w[56]), .i3(stg1_c6_w[55]), .ci(stg2_co3[63]), .s(stg2_s3[64]), .c(stg2_c3[64]), .co(stg2_co3[64]));
counter_5to3 u_a23_65(.i0(stg1_s5_w[65]), .i1(stg1_c5_w[64]), .i2(stg1_s6_w[57]), .i3(stg1_c6_w[56]), .ci(stg2_co3[64]), .s(stg2_s3[65]), .c(stg2_c3[65]), .co(stg2_co3[65]));
counter_5to3 u_a23_66(.i0(stg1_s5_w[66]), .i1(stg1_c5_w[65]), .i2(stg1_s6_w[58]), .i3(stg1_c6_w[57]), .ci(stg2_co3[65]), .s(stg2_s3[66]), .c(stg2_c3[66]), .co(stg2_co3[66]));
counter_5to3 u_a23_67(.i0(stg1_s5_w[67]), .i1(stg1_c5_w[66]), .i2(stg1_s6_w[59]), .i3(stg1_c6_w[58]), .ci(stg2_co3[66]), .s(stg2_s3[67]), .c(stg2_c3[67]), .co(stg2_co3[67]));
counter_5to3 u_a23_68(.i0(stg1_s5_w[68]), .i1(stg1_c5_w[67]), .i2(stg1_s6_w[60]), .i3(stg1_c6_w[59]), .ci(stg2_co3[67]), .s(stg2_s3[68]), .c(stg2_c3[68]), .co(stg2_co3[68]));
counter_5to3 u_a23_69(.i0(stg1_s5_w[69]), .i1(stg1_c5_w[68]), .i2(stg1_s6_w[61]), .i3(stg1_c6_w[60]), .ci(stg2_co3[68]), .s(stg2_s3[69]), .c(stg2_c3[69]), .co(stg2_co3[69]));
counter_5to3 u_a23_70(.i0(stg1_s5_w[70]), .i1(stg1_c5_w[69]), .i2(stg1_s6_w[62]), .i3(stg1_c6_w[61]), .ci(stg2_co3[69]), .s(stg2_s3[70]), .c(stg2_c3[70]), .co(stg2_co3[70]));
counter_5to3 u_a23_71(.i0(stg1_s5_w[71]), .i1(stg1_c5_w[70]), .i2(stg1_s6_w[63]), .i3(stg1_c6_w[62]), .ci(stg2_co3[70]), .s(stg2_s3[71]), .c(stg2_c3[71]), .co(stg2_co3[71]));
counter_5to3 u_a23_72(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[71]), .i2(stg1_s6_w[64]), .i3(stg1_c6_w[63]), .ci(stg2_co3[71]), .s(stg2_s3[72]), .c(stg2_c3[72]), .co(stg2_co3[72]));
counter_5to3 u_a23_73(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[65]), .i3(stg1_c6_w[64]), .ci(stg2_co3[72]), .s(stg2_s3[73]), .c(stg2_c3[73]), .co(stg2_co3[73]));
counter_5to3 u_a23_74(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[66]), .i3(stg1_c6_w[65]), .ci(stg2_co3[73]), .s(stg2_s3[74]), .c(stg2_c3[74]), .co(stg2_co3[74]));
counter_5to3 u_a23_75(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[67]), .i3(stg1_c6_w[66]), .ci(stg2_co3[74]), .s(stg2_s3[75]), .c(stg2_c3[75]), .co(stg2_co3[75]));
counter_5to3 u_a23_76(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[68]), .i3(stg1_c6_w[67]), .ci(stg2_co3[75]), .s(stg2_s3[76]), .c(stg2_c3[76]), .co(stg2_co3[76]));
counter_5to3 u_a23_77(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[69]), .i3(stg1_c6_w[68]), .ci(stg2_co3[76]), .s(stg2_s3[77]), .c(stg2_c3[77]), .co(stg2_co3[77]));
counter_5to3 u_a23_78(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[70]), .i3(stg1_c6_w[69]), .ci(stg2_co3[77]), .s(stg2_s3[78]), .c(stg2_c3[78]), .co(stg2_co3[78]));
counter_5to3 u_a23_79(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[71]), .i3(stg1_c6_w[70]), .ci(stg2_co3[78]), .s(stg2_s3[79]), .c(stg2_c3[79]), .co(stg2_co3[79]));
counter_5to3 u_a23_80(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[72]), .i3(stg1_c6_w[71]), .ci(stg2_co3[79]), .s(stg2_s3[80]), .c(stg2_c3[80]), .co(stg2_co3[80]));
counter_5to3 u_a23_81(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[72]), .i3(stg1_c6_w[72]), .ci(stg2_co3[80]), .s(stg2_s3[81]), .c(stg2_c3[81]), .co(stg2_co3[81]));
counter_5to3 u_a23_82(.i0(stg1_s5_w[72]), .i1(stg1_c5_w[72]), .i2(stg1_s6_w[72]), .i3(stg1_c6_w[72]), .ci(stg2_co3[81]), .s(stg2_s3[82]), .c(stg2_c3[82]), .co(stg2_co3[82]));

// =========================== second stage 4th group ============================================================================================================
counter_5to3 u_a24_0 (.i0(stg1_s7_w[0 ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0         ), .ci(1'b0        ), .s(stg2_s4[0 ]), .c(stg2_c4[0 ]), .co(stg2_co4[0 ]));
counter_5to3 u_a24_1 (.i0(stg1_s7_w[1 ]), .i1(stg1_c7_w[0 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[0 ]), .s(stg2_s4[1 ]), .c(stg2_c4[1 ]), .co(stg2_co4[1 ]));
counter_5to3 u_a24_2 (.i0(stg1_s7_w[2 ]), .i1(stg1_c7_w[1 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[1 ]), .s(stg2_s4[2 ]), .c(stg2_c4[2 ]), .co(stg2_co4[2 ]));
counter_5to3 u_a24_3 (.i0(stg1_s7_w[3 ]), .i1(stg1_c7_w[2 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[2 ]), .s(stg2_s4[3 ]), .c(stg2_c4[3 ]), .co(stg2_co4[3 ]));
counter_5to3 u_a24_4 (.i0(stg1_s7_w[4 ]), .i1(stg1_c7_w[3 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[3 ]), .s(stg2_s4[4 ]), .c(stg2_c4[4 ]), .co(stg2_co4[4 ]));
counter_5to3 u_a24_5 (.i0(stg1_s7_w[5 ]), .i1(stg1_c7_w[4 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[4 ]), .s(stg2_s4[5 ]), .c(stg2_c4[5 ]), .co(stg2_co4[5 ]));
counter_5to3 u_a24_6 (.i0(stg1_s7_w[6 ]), .i1(stg1_c7_w[5 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[5 ]), .s(stg2_s4[6 ]), .c(stg2_c4[6 ]), .co(stg2_co4[6 ]));
counter_5to3 u_a24_7 (.i0(stg1_s7_w[7 ]), .i1(stg1_c7_w[6 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg2_co4[6 ]), .s(stg2_s4[7 ]), .c(stg2_c4[7 ]), .co(stg2_co4[7 ]));
counter_5to3 u_a24_8 (.i0(stg1_s7_w[8 ]), .i1(stg1_c7_w[7 ]), .i2(stg1_s8_w[0 ]), .i3(1'b0         ), .ci(stg2_co4[7 ]), .s(stg2_s4[8 ]), .c(stg2_c4[8 ]), .co(stg2_co4[8 ]));
counter_5to3 u_a24_9 (.i0(stg1_s7_w[9 ]), .i1(stg1_c7_w[8 ]), .i2(stg1_s8_w[1 ]), .i3(stg1_c8_w[0 ]), .ci(stg2_co4[8 ]), .s(stg2_s4[9 ]), .c(stg2_c4[9 ]), .co(stg2_co4[9 ]));
counter_5to3 u_a24_10(.i0(stg1_s7_w[10]), .i1(stg1_c7_w[9 ]), .i2(stg1_s8_w[2 ]), .i3(stg1_c8_w[1 ]), .ci(stg2_co4[9 ]), .s(stg2_s4[10]), .c(stg2_c4[10]), .co(stg2_co4[10]));
counter_5to3 u_a24_11(.i0(stg1_s7_w[11]), .i1(stg1_c7_w[10]), .i2(stg1_s8_w[3 ]), .i3(stg1_c8_w[2 ]), .ci(stg2_co4[10]), .s(stg2_s4[11]), .c(stg2_c4[11]), .co(stg2_co4[11]));
counter_5to3 u_a24_12(.i0(stg1_s7_w[12]), .i1(stg1_c7_w[11]), .i2(stg1_s8_w[4 ]), .i3(stg1_c8_w[3 ]), .ci(stg2_co4[11]), .s(stg2_s4[12]), .c(stg2_c4[12]), .co(stg2_co4[12]));
counter_5to3 u_a24_13(.i0(stg1_s7_w[13]), .i1(stg1_c7_w[12]), .i2(stg1_s8_w[5 ]), .i3(stg1_c8_w[4 ]), .ci(stg2_co4[12]), .s(stg2_s4[13]), .c(stg2_c4[13]), .co(stg2_co4[13]));
counter_5to3 u_a24_14(.i0(stg1_s7_w[14]), .i1(stg1_c7_w[13]), .i2(stg1_s8_w[6 ]), .i3(stg1_c8_w[5 ]), .ci(stg2_co4[13]), .s(stg2_s4[14]), .c(stg2_c4[14]), .co(stg2_co4[14]));
counter_5to3 u_a24_15(.i0(stg1_s7_w[15]), .i1(stg1_c7_w[14]), .i2(stg1_s8_w[7 ]), .i3(stg1_c8_w[6 ]), .ci(stg2_co4[14]), .s(stg2_s4[15]), .c(stg2_c4[15]), .co(stg2_co4[15]));
counter_5to3 u_a24_16(.i0(stg1_s7_w[16]), .i1(stg1_c7_w[15]), .i2(stg1_s8_w[8 ]), .i3(stg1_c8_w[7 ]), .ci(stg2_co4[15]), .s(stg2_s4[16]), .c(stg2_c4[16]), .co(stg2_co4[16]));
counter_5to3 u_a24_17(.i0(stg1_s7_w[17]), .i1(stg1_c7_w[16]), .i2(stg1_s8_w[9 ]), .i3(stg1_c8_w[8 ]), .ci(stg2_co4[16]), .s(stg2_s4[17]), .c(stg2_c4[17]), .co(stg2_co4[17]));
counter_5to3 u_a24_18(.i0(stg1_s7_w[18]), .i1(stg1_c7_w[17]), .i2(stg1_s8_w[10]), .i3(stg1_c8_w[9 ]), .ci(stg2_co4[17]), .s(stg2_s4[18]), .c(stg2_c4[18]), .co(stg2_co4[18]));
counter_5to3 u_a24_19(.i0(stg1_s7_w[19]), .i1(stg1_c7_w[18]), .i2(stg1_s8_w[11]), .i3(stg1_c8_w[10]), .ci(stg2_co4[18]), .s(stg2_s4[19]), .c(stg2_c4[19]), .co(stg2_co4[19]));
counter_5to3 u_a24_20(.i0(stg1_s7_w[20]), .i1(stg1_c7_w[19]), .i2(stg1_s8_w[12]), .i3(stg1_c8_w[11]), .ci(stg2_co4[19]), .s(stg2_s4[20]), .c(stg2_c4[20]), .co(stg2_co4[20]));
counter_5to3 u_a24_21(.i0(stg1_s7_w[21]), .i1(stg1_c7_w[20]), .i2(stg1_s8_w[13]), .i3(stg1_c8_w[12]), .ci(stg2_co4[20]), .s(stg2_s4[21]), .c(stg2_c4[21]), .co(stg2_co4[21]));
counter_5to3 u_a24_22(.i0(stg1_s7_w[22]), .i1(stg1_c7_w[21]), .i2(stg1_s8_w[14]), .i3(stg1_c8_w[13]), .ci(stg2_co4[21]), .s(stg2_s4[22]), .c(stg2_c4[22]), .co(stg2_co4[22]));
counter_5to3 u_a24_23(.i0(stg1_s7_w[23]), .i1(stg1_c7_w[22]), .i2(stg1_s8_w[15]), .i3(stg1_c8_w[14]), .ci(stg2_co4[22]), .s(stg2_s4[23]), .c(stg2_c4[23]), .co(stg2_co4[23]));
counter_5to3 u_a24_24(.i0(stg1_s7_w[24]), .i1(stg1_c7_w[23]), .i2(stg1_s8_w[16]), .i3(stg1_c8_w[15]), .ci(stg2_co4[23]), .s(stg2_s4[24]), .c(stg2_c4[24]), .co(stg2_co4[24]));
counter_5to3 u_a24_25(.i0(stg1_s7_w[25]), .i1(stg1_c7_w[24]), .i2(stg1_s8_w[17]), .i3(stg1_c8_w[16]), .ci(stg2_co4[24]), .s(stg2_s4[25]), .c(stg2_c4[25]), .co(stg2_co4[25]));
counter_5to3 u_a24_26(.i0(stg1_s7_w[26]), .i1(stg1_c7_w[25]), .i2(stg1_s8_w[18]), .i3(stg1_c8_w[17]), .ci(stg2_co4[25]), .s(stg2_s4[26]), .c(stg2_c4[26]), .co(stg2_co4[26]));
counter_5to3 u_a24_27(.i0(stg1_s7_w[27]), .i1(stg1_c7_w[26]), .i2(stg1_s8_w[19]), .i3(stg1_c8_w[18]), .ci(stg2_co4[26]), .s(stg2_s4[27]), .c(stg2_c4[27]), .co(stg2_co4[27]));
counter_5to3 u_a24_28(.i0(stg1_s7_w[28]), .i1(stg1_c7_w[27]), .i2(stg1_s8_w[20]), .i3(stg1_c8_w[19]), .ci(stg2_co4[27]), .s(stg2_s4[28]), .c(stg2_c4[28]), .co(stg2_co4[28]));
counter_5to3 u_a24_29(.i0(stg1_s7_w[29]), .i1(stg1_c7_w[28]), .i2(stg1_s8_w[21]), .i3(stg1_c8_w[20]), .ci(stg2_co4[28]), .s(stg2_s4[29]), .c(stg2_c4[29]), .co(stg2_co4[29]));
counter_5to3 u_a24_30(.i0(stg1_s7_w[30]), .i1(stg1_c7_w[29]), .i2(stg1_s8_w[22]), .i3(stg1_c8_w[21]), .ci(stg2_co4[29]), .s(stg2_s4[30]), .c(stg2_c4[30]), .co(stg2_co4[30]));
counter_5to3 u_a24_31(.i0(stg1_s7_w[31]), .i1(stg1_c7_w[30]), .i2(stg1_s8_w[23]), .i3(stg1_c8_w[22]), .ci(stg2_co4[30]), .s(stg2_s4[31]), .c(stg2_c4[31]), .co(stg2_co4[31]));
counter_5to3 u_a24_32(.i0(stg1_s7_w[32]), .i1(stg1_c7_w[31]), .i2(stg1_s8_w[24]), .i3(stg1_c8_w[23]), .ci(stg2_co4[31]), .s(stg2_s4[32]), .c(stg2_c4[32]), .co(stg2_co4[32]));
counter_5to3 u_a24_33(.i0(stg1_s7_w[33]), .i1(stg1_c7_w[32]), .i2(stg1_s8_w[25]), .i3(stg1_c8_w[24]), .ci(stg2_co4[32]), .s(stg2_s4[33]), .c(stg2_c4[33]), .co(stg2_co4[33]));
counter_5to3 u_a24_34(.i0(stg1_s7_w[34]), .i1(stg1_c7_w[33]), .i2(stg1_s8_w[26]), .i3(stg1_c8_w[25]), .ci(stg2_co4[33]), .s(stg2_s4[34]), .c(stg2_c4[34]), .co(stg2_co4[34]));
counter_5to3 u_a24_35(.i0(stg1_s7_w[35]), .i1(stg1_c7_w[34]), .i2(stg1_s8_w[27]), .i3(stg1_c8_w[26]), .ci(stg2_co4[34]), .s(stg2_s4[35]), .c(stg2_c4[35]), .co(stg2_co4[35]));
counter_5to3 u_a24_36(.i0(stg1_s7_w[36]), .i1(stg1_c7_w[35]), .i2(stg1_s8_w[28]), .i3(stg1_c8_w[27]), .ci(stg2_co4[35]), .s(stg2_s4[36]), .c(stg2_c4[36]), .co(stg2_co4[36]));
counter_5to3 u_a24_37(.i0(stg1_s7_w[37]), .i1(stg1_c7_w[36]), .i2(stg1_s8_w[29]), .i3(stg1_c8_w[28]), .ci(stg2_co4[36]), .s(stg2_s4[37]), .c(stg2_c4[37]), .co(stg2_co4[37]));
counter_5to3 u_a24_38(.i0(stg1_s7_w[38]), .i1(stg1_c7_w[37]), .i2(stg1_s8_w[30]), .i3(stg1_c8_w[29]), .ci(stg2_co4[37]), .s(stg2_s4[38]), .c(stg2_c4[38]), .co(stg2_co4[38]));
counter_5to3 u_a24_39(.i0(stg1_s7_w[39]), .i1(stg1_c7_w[38]), .i2(stg1_s8_w[31]), .i3(stg1_c8_w[30]), .ci(stg2_co4[38]), .s(stg2_s4[39]), .c(stg2_c4[39]), .co(stg2_co4[39]));
counter_5to3 u_a24_40(.i0(stg1_s7_w[40]), .i1(stg1_c7_w[39]), .i2(stg1_s8_w[32]), .i3(stg1_c8_w[31]), .ci(stg2_co4[39]), .s(stg2_s4[40]), .c(stg2_c4[40]), .co(stg2_co4[40]));
counter_5to3 u_a24_41(.i0(stg1_s7_w[41]), .i1(stg1_c7_w[40]), .i2(stg1_s8_w[33]), .i3(stg1_c8_w[32]), .ci(stg2_co4[40]), .s(stg2_s4[41]), .c(stg2_c4[41]), .co(stg2_co4[41]));
counter_5to3 u_a24_42(.i0(stg1_s7_w[42]), .i1(stg1_c7_w[41]), .i2(stg1_s8_w[34]), .i3(stg1_c8_w[33]), .ci(stg2_co4[41]), .s(stg2_s4[42]), .c(stg2_c4[42]), .co(stg2_co4[42]));
counter_5to3 u_a24_43(.i0(stg1_s7_w[43]), .i1(stg1_c7_w[42]), .i2(stg1_s8_w[35]), .i3(stg1_c8_w[34]), .ci(stg2_co4[42]), .s(stg2_s4[43]), .c(stg2_c4[43]), .co(stg2_co4[43]));
counter_5to3 u_a24_44(.i0(stg1_s7_w[44]), .i1(stg1_c7_w[43]), .i2(stg1_s8_w[36]), .i3(stg1_c8_w[35]), .ci(stg2_co4[43]), .s(stg2_s4[44]), .c(stg2_c4[44]), .co(stg2_co4[44]));
counter_5to3 u_a24_45(.i0(stg1_s7_w[45]), .i1(stg1_c7_w[44]), .i2(stg1_s8_w[37]), .i3(stg1_c8_w[36]), .ci(stg2_co4[44]), .s(stg2_s4[45]), .c(stg2_c4[45]), .co(stg2_co4[45]));
counter_5to3 u_a24_46(.i0(stg1_s7_w[46]), .i1(stg1_c7_w[45]), .i2(stg1_s8_w[38]), .i3(stg1_c8_w[37]), .ci(stg2_co4[45]), .s(stg2_s4[46]), .c(stg2_c4[46]), .co(stg2_co4[46]));
counter_5to3 u_a24_47(.i0(stg1_s7_w[47]), .i1(stg1_c7_w[46]), .i2(stg1_s8_w[39]), .i3(stg1_c8_w[38]), .ci(stg2_co4[46]), .s(stg2_s4[47]), .c(stg2_c4[47]), .co(stg2_co4[47]));
counter_5to3 u_a24_48(.i0(stg1_s7_w[48]), .i1(stg1_c7_w[47]), .i2(stg1_s8_w[40]), .i3(stg1_c8_w[39]), .ci(stg2_co4[47]), .s(stg2_s4[48]), .c(stg2_c4[48]), .co(stg2_co4[48]));
counter_5to3 u_a24_49(.i0(stg1_s7_w[49]), .i1(stg1_c7_w[48]), .i2(stg1_s8_w[41]), .i3(stg1_c8_w[40]), .ci(stg2_co4[48]), .s(stg2_s4[49]), .c(stg2_c4[49]), .co(stg2_co4[49]));
counter_5to3 u_a24_50(.i0(stg1_s7_w[50]), .i1(stg1_c7_w[49]), .i2(stg1_s8_w[42]), .i3(stg1_c8_w[41]), .ci(stg2_co4[49]), .s(stg2_s4[50]), .c(stg2_c4[50]), .co(stg2_co4[50]));
counter_5to3 u_a24_51(.i0(stg1_s7_w[51]), .i1(stg1_c7_w[50]), .i2(stg1_s8_w[43]), .i3(stg1_c8_w[42]), .ci(stg2_co4[50]), .s(stg2_s4[51]), .c(stg2_c4[51]), .co(stg2_co4[51]));
counter_5to3 u_a24_52(.i0(stg1_s7_w[52]), .i1(stg1_c7_w[51]), .i2(stg1_s8_w[44]), .i3(stg1_c8_w[43]), .ci(stg2_co4[51]), .s(stg2_s4[52]), .c(stg2_c4[52]), .co(stg2_co4[52]));
counter_5to3 u_a24_53(.i0(stg1_s7_w[53]), .i1(stg1_c7_w[52]), .i2(stg1_s8_w[45]), .i3(stg1_c8_w[44]), .ci(stg2_co4[52]), .s(stg2_s4[53]), .c(stg2_c4[53]), .co(stg2_co4[53]));
counter_5to3 u_a24_54(.i0(stg1_s7_w[54]), .i1(stg1_c7_w[53]), .i2(stg1_s8_w[46]), .i3(stg1_c8_w[45]), .ci(stg2_co4[53]), .s(stg2_s4[54]), .c(stg2_c4[54]), .co(stg2_co4[54]));
counter_5to3 u_a24_55(.i0(stg1_s7_w[55]), .i1(stg1_c7_w[54]), .i2(stg1_s8_w[47]), .i3(stg1_c8_w[46]), .ci(stg2_co4[54]), .s(stg2_s4[55]), .c(stg2_c4[55]), .co(stg2_co4[55]));
counter_5to3 u_a24_56(.i0(stg1_s7_w[56]), .i1(stg1_c7_w[55]), .i2(stg1_s8_w[48]), .i3(stg1_c8_w[47]), .ci(stg2_co4[55]), .s(stg2_s4[56]), .c(stg2_c4[56]), .co(stg2_co4[56]));
counter_5to3 u_a24_57(.i0(stg1_s7_w[57]), .i1(stg1_c7_w[56]), .i2(stg1_s8_w[49]), .i3(stg1_c8_w[48]), .ci(stg2_co4[56]), .s(stg2_s4[57]), .c(stg2_c4[57]), .co(stg2_co4[57]));
counter_5to3 u_a24_58(.i0(stg1_s7_w[58]), .i1(stg1_c7_w[57]), .i2(stg1_s8_w[50]), .i3(stg1_c8_w[49]), .ci(stg2_co4[57]), .s(stg2_s4[58]), .c(stg2_c4[58]), .co(stg2_co4[58]));
counter_5to3 u_a24_59(.i0(stg1_s7_w[59]), .i1(stg1_c7_w[58]), .i2(stg1_s8_w[51]), .i3(stg1_c8_w[50]), .ci(stg2_co4[58]), .s(stg2_s4[59]), .c(stg2_c4[59]), .co(stg2_co4[59]));
counter_5to3 u_a24_60(.i0(stg1_s7_w[60]), .i1(stg1_c7_w[59]), .i2(stg1_s8_w[52]), .i3(stg1_c8_w[51]), .ci(stg2_co4[59]), .s(stg2_s4[60]), .c(stg2_c4[60]), .co(stg2_co4[60]));
counter_5to3 u_a24_61(.i0(stg1_s7_w[61]), .i1(stg1_c7_w[60]), .i2(stg1_s8_w[53]), .i3(stg1_c8_w[52]), .ci(stg2_co4[60]), .s(stg2_s4[61]), .c(stg2_c4[61]), .co(stg2_co4[61]));
counter_5to3 u_a24_62(.i0(stg1_s7_w[62]), .i1(stg1_c7_w[61]), .i2(stg1_s8_w[54]), .i3(stg1_c8_w[53]), .ci(stg2_co4[61]), .s(stg2_s4[62]), .c(stg2_c4[62]), .co(stg2_co4[62]));
counter_5to3 u_a24_63(.i0(stg1_s7_w[63]), .i1(stg1_c7_w[62]), .i2(stg1_s8_w[55]), .i3(stg1_c8_w[54]), .ci(stg2_co4[62]), .s(stg2_s4[63]), .c(stg2_c4[63]), .co(stg2_co4[63]));
counter_5to3 u_a24_64(.i0(stg1_s7_w[64]), .i1(stg1_c7_w[63]), .i2(stg1_s8_w[56]), .i3(stg1_c8_w[55]), .ci(stg2_co4[63]), .s(stg2_s4[64]), .c(stg2_c4[64]), .co(stg2_co4[64]));
counter_5to3 u_a24_65(.i0(stg1_s7_w[65]), .i1(stg1_c7_w[64]), .i2(stg1_s8_w[57]), .i3(stg1_c8_w[56]), .ci(stg2_co4[64]), .s(stg2_s4[65]), .c(stg2_c4[65]), .co(stg2_co4[65]));
counter_5to3 u_a24_66(.i0(stg1_s7_w[66]), .i1(stg1_c7_w[65]), .i2(stg1_s8_w[58]), .i3(stg1_c8_w[57]), .ci(stg2_co4[65]), .s(stg2_s4[66]), .c(stg2_c4[66]), .co(stg2_co4[66]));
counter_5to3 u_a24_67(.i0(stg1_s7_w[67]), .i1(stg1_c7_w[66]), .i2(stg1_s8_w[59]), .i3(stg1_c8_w[58]), .ci(stg2_co4[66]), .s(stg2_s4[67]), .c(stg2_c4[67]), .co(stg2_co4[67]));
counter_5to3 u_a24_68(.i0(stg1_s7_w[68]), .i1(stg1_c7_w[67]), .i2(stg1_s8_w[60]), .i3(stg1_c8_w[59]), .ci(stg2_co4[67]), .s(stg2_s4[68]), .c(stg2_c4[68]), .co(stg2_co4[68]));
counter_5to3 u_a24_69(.i0(stg1_s7_w[69]), .i1(stg1_c7_w[68]), .i2(stg1_s8_w[61]), .i3(stg1_c8_w[60]), .ci(stg2_co4[68]), .s(stg2_s4[69]), .c(stg2_c4[69]), .co(stg2_co4[69]));
counter_5to3 u_a24_70(.i0(stg1_s7_w[70]), .i1(stg1_c7_w[69]), .i2(stg1_s8_w[62]), .i3(stg1_c8_w[61]), .ci(stg2_co4[69]), .s(stg2_s4[70]), .c(stg2_c4[70]), .co(stg2_co4[70]));
counter_5to3 u_a24_71(.i0(stg1_s7_w[71]), .i1(stg1_c7_w[70]), .i2(stg1_s8_w[63]), .i3(stg1_c8_w[62]), .ci(stg2_co4[70]), .s(stg2_s4[71]), .c(stg2_c4[71]), .co(stg2_co4[71]));
counter_5to3 u_a24_72(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[71]), .i2(stg1_s8_w[64]), .i3(stg1_c8_w[63]), .ci(stg2_co4[71]), .s(stg2_s4[72]), .c(stg2_c4[72]), .co(stg2_co4[72]));
counter_5to3 u_a24_73(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[65]), .i3(stg1_c8_w[64]), .ci(stg2_co4[72]), .s(stg2_s4[73]), .c(stg2_c4[73]), .co(stg2_co4[73]));
counter_5to3 u_a24_74(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[66]), .i3(stg1_c8_w[65]), .ci(stg2_co4[73]), .s(stg2_s4[74]), .c(stg2_c4[74]), .co(stg2_co4[74]));
counter_5to3 u_a24_75(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[67]), .i3(stg1_c8_w[66]), .ci(stg2_co4[74]), .s(stg2_s4[75]), .c(stg2_c4[75]), .co(stg2_co4[75]));
counter_5to3 u_a24_76(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[68]), .i3(stg1_c8_w[67]), .ci(stg2_co4[75]), .s(stg2_s4[76]), .c(stg2_c4[76]), .co(stg2_co4[76]));
counter_5to3 u_a24_77(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[69]), .i3(stg1_c8_w[68]), .ci(stg2_co4[76]), .s(stg2_s4[77]), .c(stg2_c4[77]), .co(stg2_co4[77]));
counter_5to3 u_a24_78(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[70]), .i3(stg1_c8_w[69]), .ci(stg2_co4[77]), .s(stg2_s4[78]), .c(stg2_c4[78]), .co(stg2_co4[78]));
counter_5to3 u_a24_79(.i0(stg1_s7_w[72]), .i1(stg1_c7_w[72]), .i2(stg1_s8_w[71]), .i3(stg1_c8_w[70]), .ci(stg2_co4[78]), .s(stg2_s4[79]), .c(stg2_c4[79]), .co(stg2_co4[79]));

//================ third stage ================
wire [82:0] stg2_s1_w, stg2_c1_w;
wire [82:0] stg2_s2_w, stg2_c2_w;
wire [82:0] stg2_s3_w, stg2_c3_w;
wire [79:0] stg2_s4_w, stg2_c4_w;
wire [65:0] pp33_w2;

// ==========pipeline ================
reg [82:0] stg2_s1_ff, stg2_c1_ff;
reg [82:0] stg2_s2_ff, stg2_c2_ff;
reg [82:0] stg2_s3_ff, stg2_c3_ff;
reg [79:0] stg2_s4_ff, stg2_c4_ff;
reg [65:0] pp33_f2;

always @(posedge clk or negedge rstn)begin
    if (!rstn)begin
        stg2_s1_ff <= 83'b0;
        stg2_c1_ff <= 83'b0;
        stg2_s2_ff <= 83'b0;
        stg2_c2_ff <= 83'b0;
        stg2_s3_ff <= 83'b0;
        stg2_c3_ff <= 83'b0;
        stg2_s4_ff <= 80'b0;
        stg2_c4_ff <= 80'b0;
        pp33_f2    <= 66'b0;
    end
    else begin
        stg2_s1_ff <= stg2_s1;
        stg2_c1_ff <= stg2_c1;
        stg2_s2_ff <= stg2_s2;
        stg2_c2_ff <= stg2_c2;
        stg2_s3_ff <= stg2_s3;
        stg2_c3_ff <= stg2_c3;
        stg2_s4_ff <= stg2_s4;
        stg2_c4_ff <= stg2_c4;
        pp33_f2    <= pp33_w1;
    end
end

assign stg2_s1_w   = stg2_s1_ff;
assign stg2_c1_w   = stg2_c1_ff;
assign stg2_s2_w   = stg2_s2_ff;
assign stg2_c2_w   = stg2_c2_ff;
assign stg2_s3_w   = stg2_s3_ff;
assign stg2_c3_w   = stg2_c3_ff;
assign stg2_s4_w   = stg2_s4_ff;
assign stg2_c4_w   = stg2_c4_ff;
assign pp33_w2     = pp33_f2   ;

wire [100:0] stg3_s1, stg3_c1, stg3_co1;
wire  [95:0] stg3_s2, stg3_c2, stg3_co2;

// =========================== third stage 1st group ============================================================================================================
counter_5to3 u_a31_0  (.i0(stg2_s1_w[0 ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0         ), .ci(1'b0        ), .s(stg3_s1[0  ]), .c(stg3_c1[0  ]), .co(stg3_co1[0  ]));
counter_5to3 u_a31_1  (.i0(stg2_s1_w[1 ]), .i1(stg2_c1_w[0 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[0 ]), .s(stg3_s1[1  ]), .c(stg3_c1[1  ]), .co(stg3_co1[1  ]));
counter_5to3 u_a31_2  (.i0(stg2_s1_w[2 ]), .i1(stg2_c1_w[1 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[1 ]), .s(stg3_s1[2  ]), .c(stg3_c1[2  ]), .co(stg3_co1[2  ]));
counter_5to3 u_a31_3  (.i0(stg2_s1_w[3 ]), .i1(stg2_c1_w[2 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[2 ]), .s(stg3_s1[3  ]), .c(stg3_c1[3  ]), .co(stg3_co1[3  ]));
counter_5to3 u_a31_4  (.i0(stg2_s1_w[4 ]), .i1(stg2_c1_w[3 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[3 ]), .s(stg3_s1[4  ]), .c(stg3_c1[4  ]), .co(stg3_co1[4  ]));
counter_5to3 u_a31_5  (.i0(stg2_s1_w[5 ]), .i1(stg2_c1_w[4 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[4 ]), .s(stg3_s1[5  ]), .c(stg3_c1[5  ]), .co(stg3_co1[5  ]));
counter_5to3 u_a31_6  (.i0(stg2_s1_w[6 ]), .i1(stg2_c1_w[5 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[5 ]), .s(stg3_s1[6  ]), .c(stg3_c1[6  ]), .co(stg3_co1[6  ]));
counter_5to3 u_a31_7  (.i0(stg2_s1_w[7 ]), .i1(stg2_c1_w[6 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[6 ]), .s(stg3_s1[7  ]), .c(stg3_c1[7  ]), .co(stg3_co1[7  ]));
counter_5to3 u_a31_8  (.i0(stg2_s1_w[8 ]), .i1(stg2_c1_w[7 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[7 ]), .s(stg3_s1[8  ]), .c(stg3_c1[8  ]), .co(stg3_co1[8  ]));
counter_5to3 u_a31_9  (.i0(stg2_s1_w[9 ]), .i1(stg2_c1_w[8 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[8 ]), .s(stg3_s1[9  ]), .c(stg3_c1[9  ]), .co(stg3_co1[9  ]));
counter_5to3 u_a31_10 (.i0(stg2_s1_w[10]), .i1(stg2_c1_w[9 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[9 ]), .s(stg3_s1[10 ]), .c(stg3_c1[10 ]), .co(stg3_co1[10 ]));
counter_5to3 u_a31_11 (.i0(stg2_s1_w[11]), .i1(stg2_c1_w[10]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[10]), .s(stg3_s1[11 ]), .c(stg3_c1[11 ]), .co(stg3_co1[11 ]));
counter_5to3 u_a31_12 (.i0(stg2_s1_w[12]), .i1(stg2_c1_w[11]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[11]), .s(stg3_s1[12 ]), .c(stg3_c1[12 ]), .co(stg3_co1[12 ]));
counter_5to3 u_a31_13 (.i0(stg2_s1_w[13]), .i1(stg2_c1_w[12]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[12]), .s(stg3_s1[13 ]), .c(stg3_c1[13 ]), .co(stg3_co1[13 ]));
counter_5to3 u_a31_14 (.i0(stg2_s1_w[14]), .i1(stg2_c1_w[13]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[13]), .s(stg3_s1[14 ]), .c(stg3_c1[14 ]), .co(stg3_co1[14 ]));
counter_5to3 u_a31_15 (.i0(stg2_s1_w[15]), .i1(stg2_c1_w[14]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co1[14]), .s(stg3_s1[15 ]), .c(stg3_c1[15 ]), .co(stg3_co1[15 ]));
counter_5to3 u_a31_16 (.i0(stg2_s1_w[16]), .i1(stg2_c1_w[15]), .i2(stg2_s2_w[0 ]), .i3(1'b0         ), .ci(stg3_co1[15]), .s(stg3_s1[16 ]), .c(stg3_c1[16 ]), .co(stg3_co1[16 ]));
counter_5to3 u_a31_17 (.i0(stg2_s1_w[17]), .i1(stg2_c1_w[16]), .i2(stg2_s2_w[1 ]), .i3(stg2_c2_w[0 ]), .ci(stg3_co1[16]), .s(stg3_s1[17 ]), .c(stg3_c1[17 ]), .co(stg3_co1[17 ]));
counter_5to3 u_a31_18 (.i0(stg2_s1_w[18]), .i1(stg2_c1_w[17]), .i2(stg2_s2_w[2 ]), .i3(stg2_c2_w[1 ]), .ci(stg3_co1[17]), .s(stg3_s1[18 ]), .c(stg3_c1[18 ]), .co(stg3_co1[18 ]));
counter_5to3 u_a31_19 (.i0(stg2_s1_w[19]), .i1(stg2_c1_w[18]), .i2(stg2_s2_w[3 ]), .i3(stg2_c2_w[2 ]), .ci(stg3_co1[18]), .s(stg3_s1[19 ]), .c(stg3_c1[19 ]), .co(stg3_co1[19 ]));
counter_5to3 u_a31_20 (.i0(stg2_s1_w[20]), .i1(stg2_c1_w[19]), .i2(stg2_s2_w[4 ]), .i3(stg2_c2_w[3 ]), .ci(stg3_co1[19]), .s(stg3_s1[20 ]), .c(stg3_c1[20 ]), .co(stg3_co1[20 ]));
counter_5to3 u_a31_21 (.i0(stg2_s1_w[21]), .i1(stg2_c1_w[20]), .i2(stg2_s2_w[5 ]), .i3(stg2_c2_w[4 ]), .ci(stg3_co1[20]), .s(stg3_s1[21 ]), .c(stg3_c1[21 ]), .co(stg3_co1[21 ]));
counter_5to3 u_a31_22 (.i0(stg2_s1_w[22]), .i1(stg2_c1_w[21]), .i2(stg2_s2_w[6 ]), .i3(stg2_c2_w[5 ]), .ci(stg3_co1[21]), .s(stg3_s1[22 ]), .c(stg3_c1[22 ]), .co(stg3_co1[22 ]));
counter_5to3 u_a31_23 (.i0(stg2_s1_w[23]), .i1(stg2_c1_w[22]), .i2(stg2_s2_w[7 ]), .i3(stg2_c2_w[6 ]), .ci(stg3_co1[22]), .s(stg3_s1[23 ]), .c(stg3_c1[23 ]), .co(stg3_co1[23 ]));
counter_5to3 u_a31_24 (.i0(stg2_s1_w[24]), .i1(stg2_c1_w[23]), .i2(stg2_s2_w[8 ]), .i3(stg2_c2_w[7 ]), .ci(stg3_co1[23]), .s(stg3_s1[24 ]), .c(stg3_c1[24 ]), .co(stg3_co1[24 ]));
counter_5to3 u_a31_25 (.i0(stg2_s1_w[25]), .i1(stg2_c1_w[24]), .i2(stg2_s2_w[9 ]), .i3(stg2_c2_w[8 ]), .ci(stg3_co1[24]), .s(stg3_s1[25 ]), .c(stg3_c1[25 ]), .co(stg3_co1[25 ]));
counter_5to3 u_a31_26 (.i0(stg2_s1_w[26]), .i1(stg2_c1_w[25]), .i2(stg2_s2_w[10]), .i3(stg2_c2_w[9 ]), .ci(stg3_co1[25]), .s(stg3_s1[26 ]), .c(stg3_c1[26 ]), .co(stg3_co1[26 ]));
counter_5to3 u_a31_27 (.i0(stg2_s1_w[27]), .i1(stg2_c1_w[26]), .i2(stg2_s2_w[11]), .i3(stg2_c2_w[10]), .ci(stg3_co1[26]), .s(stg3_s1[27 ]), .c(stg3_c1[27 ]), .co(stg3_co1[27 ]));
counter_5to3 u_a31_28 (.i0(stg2_s1_w[28]), .i1(stg2_c1_w[27]), .i2(stg2_s2_w[12]), .i3(stg2_c2_w[11]), .ci(stg3_co1[27]), .s(stg3_s1[28 ]), .c(stg3_c1[28 ]), .co(stg3_co1[28 ]));
counter_5to3 u_a31_29 (.i0(stg2_s1_w[29]), .i1(stg2_c1_w[28]), .i2(stg2_s2_w[13]), .i3(stg2_c2_w[12]), .ci(stg3_co1[28]), .s(stg3_s1[29 ]), .c(stg3_c1[29 ]), .co(stg3_co1[29 ]));
counter_5to3 u_a31_30 (.i0(stg2_s1_w[30]), .i1(stg2_c1_w[29]), .i2(stg2_s2_w[14]), .i3(stg2_c2_w[13]), .ci(stg3_co1[29]), .s(stg3_s1[30 ]), .c(stg3_c1[30 ]), .co(stg3_co1[30 ]));
counter_5to3 u_a31_31 (.i0(stg2_s1_w[31]), .i1(stg2_c1_w[30]), .i2(stg2_s2_w[15]), .i3(stg2_c2_w[14]), .ci(stg3_co1[30]), .s(stg3_s1[31 ]), .c(stg3_c1[31 ]), .co(stg3_co1[31 ]));
counter_5to3 u_a31_32 (.i0(stg2_s1_w[32]), .i1(stg2_c1_w[31]), .i2(stg2_s2_w[16]), .i3(stg2_c2_w[15]), .ci(stg3_co1[31]), .s(stg3_s1[32 ]), .c(stg3_c1[32 ]), .co(stg3_co1[32 ]));
counter_5to3 u_a31_33 (.i0(stg2_s1_w[33]), .i1(stg2_c1_w[32]), .i2(stg2_s2_w[17]), .i3(stg2_c2_w[16]), .ci(stg3_co1[32]), .s(stg3_s1[33 ]), .c(stg3_c1[33 ]), .co(stg3_co1[33 ]));
counter_5to3 u_a31_34 (.i0(stg2_s1_w[34]), .i1(stg2_c1_w[33]), .i2(stg2_s2_w[18]), .i3(stg2_c2_w[17]), .ci(stg3_co1[33]), .s(stg3_s1[34 ]), .c(stg3_c1[34 ]), .co(stg3_co1[34 ]));
counter_5to3 u_a31_35 (.i0(stg2_s1_w[35]), .i1(stg2_c1_w[34]), .i2(stg2_s2_w[19]), .i3(stg2_c2_w[18]), .ci(stg3_co1[34]), .s(stg3_s1[35 ]), .c(stg3_c1[35 ]), .co(stg3_co1[35 ]));
counter_5to3 u_a31_36 (.i0(stg2_s1_w[36]), .i1(stg2_c1_w[35]), .i2(stg2_s2_w[20]), .i3(stg2_c2_w[19]), .ci(stg3_co1[35]), .s(stg3_s1[36 ]), .c(stg3_c1[36 ]), .co(stg3_co1[36 ]));
counter_5to3 u_a31_37 (.i0(stg2_s1_w[37]), .i1(stg2_c1_w[36]), .i2(stg2_s2_w[21]), .i3(stg2_c2_w[20]), .ci(stg3_co1[36]), .s(stg3_s1[37 ]), .c(stg3_c1[37 ]), .co(stg3_co1[37 ]));
counter_5to3 u_a31_38 (.i0(stg2_s1_w[38]), .i1(stg2_c1_w[37]), .i2(stg2_s2_w[22]), .i3(stg2_c2_w[21]), .ci(stg3_co1[37]), .s(stg3_s1[38 ]), .c(stg3_c1[38 ]), .co(stg3_co1[38 ]));
counter_5to3 u_a31_39 (.i0(stg2_s1_w[39]), .i1(stg2_c1_w[38]), .i2(stg2_s2_w[23]), .i3(stg2_c2_w[22]), .ci(stg3_co1[38]), .s(stg3_s1[39 ]), .c(stg3_c1[39 ]), .co(stg3_co1[39 ]));
counter_5to3 u_a31_40 (.i0(stg2_s1_w[40]), .i1(stg2_c1_w[39]), .i2(stg2_s2_w[24]), .i3(stg2_c2_w[23]), .ci(stg3_co1[39]), .s(stg3_s1[40 ]), .c(stg3_c1[40 ]), .co(stg3_co1[40 ]));
counter_5to3 u_a31_41 (.i0(stg2_s1_w[41]), .i1(stg2_c1_w[40]), .i2(stg2_s2_w[25]), .i3(stg2_c2_w[24]), .ci(stg3_co1[40]), .s(stg3_s1[41 ]), .c(stg3_c1[41 ]), .co(stg3_co1[41 ]));
counter_5to3 u_a31_42 (.i0(stg2_s1_w[42]), .i1(stg2_c1_w[41]), .i2(stg2_s2_w[26]), .i3(stg2_c2_w[25]), .ci(stg3_co1[41]), .s(stg3_s1[42 ]), .c(stg3_c1[42 ]), .co(stg3_co1[42 ]));
counter_5to3 u_a31_43 (.i0(stg2_s1_w[43]), .i1(stg2_c1_w[42]), .i2(stg2_s2_w[27]), .i3(stg2_c2_w[26]), .ci(stg3_co1[42]), .s(stg3_s1[43 ]), .c(stg3_c1[43 ]), .co(stg3_co1[43 ]));
counter_5to3 u_a31_44 (.i0(stg2_s1_w[44]), .i1(stg2_c1_w[43]), .i2(stg2_s2_w[28]), .i3(stg2_c2_w[27]), .ci(stg3_co1[43]), .s(stg3_s1[44 ]), .c(stg3_c1[44 ]), .co(stg3_co1[44 ]));
counter_5to3 u_a31_45 (.i0(stg2_s1_w[45]), .i1(stg2_c1_w[44]), .i2(stg2_s2_w[29]), .i3(stg2_c2_w[28]), .ci(stg3_co1[44]), .s(stg3_s1[45 ]), .c(stg3_c1[45 ]), .co(stg3_co1[45 ]));
counter_5to3 u_a31_46 (.i0(stg2_s1_w[46]), .i1(stg2_c1_w[45]), .i2(stg2_s2_w[30]), .i3(stg2_c2_w[29]), .ci(stg3_co1[45]), .s(stg3_s1[46 ]), .c(stg3_c1[46 ]), .co(stg3_co1[46 ]));
counter_5to3 u_a31_47 (.i0(stg2_s1_w[47]), .i1(stg2_c1_w[46]), .i2(stg2_s2_w[31]), .i3(stg2_c2_w[30]), .ci(stg3_co1[46]), .s(stg3_s1[47 ]), .c(stg3_c1[47 ]), .co(stg3_co1[47 ]));
counter_5to3 u_a31_48 (.i0(stg2_s1_w[48]), .i1(stg2_c1_w[47]), .i2(stg2_s2_w[32]), .i3(stg2_c2_w[31]), .ci(stg3_co1[47]), .s(stg3_s1[48 ]), .c(stg3_c1[48 ]), .co(stg3_co1[48 ]));
counter_5to3 u_a31_49 (.i0(stg2_s1_w[49]), .i1(stg2_c1_w[48]), .i2(stg2_s2_w[33]), .i3(stg2_c2_w[32]), .ci(stg3_co1[48]), .s(stg3_s1[49 ]), .c(stg3_c1[49 ]), .co(stg3_co1[49 ]));
counter_5to3 u_a31_50 (.i0(stg2_s1_w[50]), .i1(stg2_c1_w[49]), .i2(stg2_s2_w[34]), .i3(stg2_c2_w[33]), .ci(stg3_co1[49]), .s(stg3_s1[50 ]), .c(stg3_c1[50 ]), .co(stg3_co1[50 ]));
counter_5to3 u_a31_51 (.i0(stg2_s1_w[51]), .i1(stg2_c1_w[50]), .i2(stg2_s2_w[35]), .i3(stg2_c2_w[34]), .ci(stg3_co1[50]), .s(stg3_s1[51 ]), .c(stg3_c1[51 ]), .co(stg3_co1[51 ]));
counter_5to3 u_a31_52 (.i0(stg2_s1_w[52]), .i1(stg2_c1_w[51]), .i2(stg2_s2_w[36]), .i3(stg2_c2_w[35]), .ci(stg3_co1[51]), .s(stg3_s1[52 ]), .c(stg3_c1[52 ]), .co(stg3_co1[52 ]));
counter_5to3 u_a31_53 (.i0(stg2_s1_w[53]), .i1(stg2_c1_w[52]), .i2(stg2_s2_w[37]), .i3(stg2_c2_w[36]), .ci(stg3_co1[52]), .s(stg3_s1[53 ]), .c(stg3_c1[53 ]), .co(stg3_co1[53 ]));
counter_5to3 u_a31_54 (.i0(stg2_s1_w[54]), .i1(stg2_c1_w[53]), .i2(stg2_s2_w[38]), .i3(stg2_c2_w[37]), .ci(stg3_co1[53]), .s(stg3_s1[54 ]), .c(stg3_c1[54 ]), .co(stg3_co1[54 ]));
counter_5to3 u_a31_55 (.i0(stg2_s1_w[55]), .i1(stg2_c1_w[54]), .i2(stg2_s2_w[39]), .i3(stg2_c2_w[38]), .ci(stg3_co1[54]), .s(stg3_s1[55 ]), .c(stg3_c1[55 ]), .co(stg3_co1[55 ]));
counter_5to3 u_a31_56 (.i0(stg2_s1_w[56]), .i1(stg2_c1_w[55]), .i2(stg2_s2_w[40]), .i3(stg2_c2_w[39]), .ci(stg3_co1[55]), .s(stg3_s1[56 ]), .c(stg3_c1[56 ]), .co(stg3_co1[56 ]));
counter_5to3 u_a31_57 (.i0(stg2_s1_w[57]), .i1(stg2_c1_w[56]), .i2(stg2_s2_w[41]), .i3(stg2_c2_w[40]), .ci(stg3_co1[56]), .s(stg3_s1[57 ]), .c(stg3_c1[57 ]), .co(stg3_co1[57 ]));
counter_5to3 u_a31_58 (.i0(stg2_s1_w[58]), .i1(stg2_c1_w[57]), .i2(stg2_s2_w[42]), .i3(stg2_c2_w[41]), .ci(stg3_co1[57]), .s(stg3_s1[58 ]), .c(stg3_c1[58 ]), .co(stg3_co1[58 ]));
counter_5to3 u_a31_59 (.i0(stg2_s1_w[59]), .i1(stg2_c1_w[58]), .i2(stg2_s2_w[43]), .i3(stg2_c2_w[42]), .ci(stg3_co1[58]), .s(stg3_s1[59 ]), .c(stg3_c1[59 ]), .co(stg3_co1[59 ]));
counter_5to3 u_a31_60 (.i0(stg2_s1_w[60]), .i1(stg2_c1_w[59]), .i2(stg2_s2_w[44]), .i3(stg2_c2_w[43]), .ci(stg3_co1[59]), .s(stg3_s1[60 ]), .c(stg3_c1[60 ]), .co(stg3_co1[60 ]));
counter_5to3 u_a31_61 (.i0(stg2_s1_w[61]), .i1(stg2_c1_w[60]), .i2(stg2_s2_w[45]), .i3(stg2_c2_w[44]), .ci(stg3_co1[60]), .s(stg3_s1[61 ]), .c(stg3_c1[61 ]), .co(stg3_co1[61 ]));
counter_5to3 u_a31_62 (.i0(stg2_s1_w[62]), .i1(stg2_c1_w[61]), .i2(stg2_s2_w[46]), .i3(stg2_c2_w[45]), .ci(stg3_co1[61]), .s(stg3_s1[62 ]), .c(stg3_c1[62 ]), .co(stg3_co1[62 ]));
counter_5to3 u_a31_63 (.i0(stg2_s1_w[63]), .i1(stg2_c1_w[62]), .i2(stg2_s2_w[47]), .i3(stg2_c2_w[46]), .ci(stg3_co1[62]), .s(stg3_s1[63 ]), .c(stg3_c1[63 ]), .co(stg3_co1[63 ]));
counter_5to3 u_a31_64 (.i0(stg2_s1_w[64]), .i1(stg2_c1_w[63]), .i2(stg2_s2_w[48]), .i3(stg2_c2_w[47]), .ci(stg3_co1[63]), .s(stg3_s1[64 ]), .c(stg3_c1[64 ]), .co(stg3_co1[64 ]));
counter_5to3 u_a31_65 (.i0(stg2_s1_w[65]), .i1(stg2_c1_w[64]), .i2(stg2_s2_w[49]), .i3(stg2_c2_w[48]), .ci(stg3_co1[64]), .s(stg3_s1[65 ]), .c(stg3_c1[65 ]), .co(stg3_co1[65 ]));
counter_5to3 u_a31_66 (.i0(stg2_s1_w[66]), .i1(stg2_c1_w[65]), .i2(stg2_s2_w[50]), .i3(stg2_c2_w[49]), .ci(stg3_co1[65]), .s(stg3_s1[66 ]), .c(stg3_c1[66 ]), .co(stg3_co1[66 ]));
counter_5to3 u_a31_67 (.i0(stg2_s1_w[67]), .i1(stg2_c1_w[66]), .i2(stg2_s2_w[51]), .i3(stg2_c2_w[50]), .ci(stg3_co1[66]), .s(stg3_s1[67 ]), .c(stg3_c1[67 ]), .co(stg3_co1[67 ]));
counter_5to3 u_a31_68 (.i0(stg2_s1_w[68]), .i1(stg2_c1_w[67]), .i2(stg2_s2_w[52]), .i3(stg2_c2_w[51]), .ci(stg3_co1[67]), .s(stg3_s1[68 ]), .c(stg3_c1[68 ]), .co(stg3_co1[68 ]));
counter_5to3 u_a31_69 (.i0(stg2_s1_w[69]), .i1(stg2_c1_w[68]), .i2(stg2_s2_w[53]), .i3(stg2_c2_w[52]), .ci(stg3_co1[68]), .s(stg3_s1[69 ]), .c(stg3_c1[69 ]), .co(stg3_co1[69 ]));
counter_5to3 u_a31_70 (.i0(stg2_s1_w[70]), .i1(stg2_c1_w[69]), .i2(stg2_s2_w[54]), .i3(stg2_c2_w[53]), .ci(stg3_co1[69]), .s(stg3_s1[70 ]), .c(stg3_c1[70 ]), .co(stg3_co1[70 ]));
counter_5to3 u_a31_71 (.i0(stg2_s1_w[71]), .i1(stg2_c1_w[70]), .i2(stg2_s2_w[55]), .i3(stg2_c2_w[54]), .ci(stg3_co1[70]), .s(stg3_s1[71 ]), .c(stg3_c1[71 ]), .co(stg3_co1[71 ]));
counter_5to3 u_a31_72 (.i0(stg2_s1_w[72]), .i1(stg2_c1_w[71]), .i2(stg2_s2_w[56]), .i3(stg2_c2_w[55]), .ci(stg3_co1[71]), .s(stg3_s1[72 ]), .c(stg3_c1[72 ]), .co(stg3_co1[72 ]));
counter_5to3 u_a31_73 (.i0(stg2_s1_w[73]), .i1(stg2_c1_w[72]), .i2(stg2_s2_w[57]), .i3(stg2_c2_w[56]), .ci(stg3_co1[72]), .s(stg3_s1[73 ]), .c(stg3_c1[73 ]), .co(stg3_co1[73 ]));
counter_5to3 u_a31_74 (.i0(stg2_s1_w[74]), .i1(stg2_c1_w[73]), .i2(stg2_s2_w[58]), .i3(stg2_c2_w[57]), .ci(stg3_co1[73]), .s(stg3_s1[74 ]), .c(stg3_c1[74 ]), .co(stg3_co1[74 ]));
counter_5to3 u_a31_75 (.i0(stg2_s1_w[75]), .i1(stg2_c1_w[74]), .i2(stg2_s2_w[59]), .i3(stg2_c2_w[58]), .ci(stg3_co1[74]), .s(stg3_s1[75 ]), .c(stg3_c1[75 ]), .co(stg3_co1[75 ]));
counter_5to3 u_a31_76 (.i0(stg2_s1_w[76]), .i1(stg2_c1_w[75]), .i2(stg2_s2_w[60]), .i3(stg2_c2_w[59]), .ci(stg3_co1[75]), .s(stg3_s1[76 ]), .c(stg3_c1[76 ]), .co(stg3_co1[76 ]));
counter_5to3 u_a31_77 (.i0(stg2_s1_w[77]), .i1(stg2_c1_w[76]), .i2(stg2_s2_w[61]), .i3(stg2_c2_w[60]), .ci(stg3_co1[76]), .s(stg3_s1[77 ]), .c(stg3_c1[77 ]), .co(stg3_co1[77 ]));
counter_5to3 u_a31_78 (.i0(stg2_s1_w[78]), .i1(stg2_c1_w[77]), .i2(stg2_s2_w[62]), .i3(stg2_c2_w[61]), .ci(stg3_co1[77]), .s(stg3_s1[78 ]), .c(stg3_c1[78 ]), .co(stg3_co1[78 ]));
counter_5to3 u_a31_79 (.i0(stg2_s1_w[79]), .i1(stg2_c1_w[78]), .i2(stg2_s2_w[63]), .i3(stg2_c2_w[62]), .ci(stg3_co1[78]), .s(stg3_s1[79 ]), .c(stg3_c1[79 ]), .co(stg3_co1[79 ]));
counter_5to3 u_a31_80 (.i0(stg2_s1_w[80]), .i1(stg2_c1_w[79]), .i2(stg2_s2_w[64]), .i3(stg2_c2_w[63]), .ci(stg3_co1[79]), .s(stg3_s1[80 ]), .c(stg3_c1[80 ]), .co(stg3_co1[80 ]));
counter_5to3 u_a31_81 (.i0(stg2_s1_w[81]), .i1(stg2_c1_w[80]), .i2(stg2_s2_w[65]), .i3(stg2_c2_w[64]), .ci(stg3_co1[80]), .s(stg3_s1[81 ]), .c(stg3_c1[81 ]), .co(stg3_co1[81 ]));
counter_5to3 u_a31_82 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[81]), .i2(stg2_s2_w[66]), .i3(stg2_c2_w[65]), .ci(stg3_co1[81]), .s(stg3_s1[82 ]), .c(stg3_c1[82 ]), .co(stg3_co1[82 ]));
counter_5to3 u_a31_83 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[67]), .i3(stg2_c2_w[66]), .ci(stg3_co1[82]), .s(stg3_s1[83 ]), .c(stg3_c1[83 ]), .co(stg3_co1[83 ]));
counter_5to3 u_a31_84 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[68]), .i3(stg2_c2_w[67]), .ci(stg3_co1[83]), .s(stg3_s1[84 ]), .c(stg3_c1[84 ]), .co(stg3_co1[84 ]));
counter_5to3 u_a31_85 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[69]), .i3(stg2_c2_w[68]), .ci(stg3_co1[84]), .s(stg3_s1[85 ]), .c(stg3_c1[85 ]), .co(stg3_co1[85 ]));
counter_5to3 u_a31_86 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[70]), .i3(stg2_c2_w[69]), .ci(stg3_co1[85]), .s(stg3_s1[86 ]), .c(stg3_c1[86 ]), .co(stg3_co1[86 ]));
counter_5to3 u_a31_87 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[71]), .i3(stg2_c2_w[70]), .ci(stg3_co1[86]), .s(stg3_s1[87 ]), .c(stg3_c1[87 ]), .co(stg3_co1[87 ]));
counter_5to3 u_a31_88 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[72]), .i3(stg2_c2_w[71]), .ci(stg3_co1[87]), .s(stg3_s1[88 ]), .c(stg3_c1[88 ]), .co(stg3_co1[88 ]));
counter_5to3 u_a31_89 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[73]), .i3(stg2_c2_w[72]), .ci(stg3_co1[88]), .s(stg3_s1[89 ]), .c(stg3_c1[89 ]), .co(stg3_co1[89 ]));
counter_5to3 u_a31_90 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[74]), .i3(stg2_c2_w[73]), .ci(stg3_co1[89]), .s(stg3_s1[90 ]), .c(stg3_c1[90 ]), .co(stg3_co1[90 ]));
counter_5to3 u_a31_91 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[75]), .i3(stg2_c2_w[74]), .ci(stg3_co1[90]), .s(stg3_s1[91 ]), .c(stg3_c1[91 ]), .co(stg3_co1[91 ]));
counter_5to3 u_a31_92 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[76]), .i3(stg2_c2_w[75]), .ci(stg3_co1[91]), .s(stg3_s1[92 ]), .c(stg3_c1[92 ]), .co(stg3_co1[92 ]));
counter_5to3 u_a31_93 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[77]), .i3(stg2_c2_w[76]), .ci(stg3_co1[92]), .s(stg3_s1[93 ]), .c(stg3_c1[93 ]), .co(stg3_co1[93 ]));
counter_5to3 u_a31_94 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[78]), .i3(stg2_c2_w[77]), .ci(stg3_co1[93]), .s(stg3_s1[94 ]), .c(stg3_c1[94 ]), .co(stg3_co1[94 ]));
counter_5to3 u_a31_95 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[79]), .i3(stg2_c2_w[78]), .ci(stg3_co1[94]), .s(stg3_s1[95 ]), .c(stg3_c1[95 ]), .co(stg3_co1[95 ]));
counter_5to3 u_a31_96 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[80]), .i3(stg2_c2_w[79]), .ci(stg3_co1[95]), .s(stg3_s1[96 ]), .c(stg3_c1[96 ]), .co(stg3_co1[96 ]));
counter_5to3 u_a31_97 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[81]), .i3(stg2_c2_w[80]), .ci(stg3_co1[96]), .s(stg3_s1[97 ]), .c(stg3_c1[97 ]), .co(stg3_co1[97 ]));
counter_5to3 u_a31_98 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[82]), .i3(stg2_c2_w[81]), .ci(stg3_co1[97]), .s(stg3_s1[98 ]), .c(stg3_c1[98 ]), .co(stg3_co1[98 ]));
counter_5to3 u_a31_99 (.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[82]), .i3(stg2_c2_w[82]), .ci(stg3_co1[98]), .s(stg3_s1[99 ]), .c(stg3_c1[99 ]), .co(stg3_co1[99 ]));
counter_5to3 u_a31_100(.i0(stg2_s1_w[82]), .i1(stg2_c1_w[82]), .i2(stg2_s2_w[82]), .i3(stg2_c2_w[82]), .ci(stg3_co1[99]), .s(stg3_s1[100]), .c(stg3_c1[100]), .co(stg3_co1[100]));

// =========================== third stage 2nd group ============================================================================================================
counter_5to3 u_a32_0  (.i0(stg2_s3_w[0 ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0         ), .ci(1'b0        ), .s(stg3_s2[0  ]), .c(stg3_c2[0  ]), .co(stg3_co2[0  ]));
counter_5to3 u_a32_1  (.i0(stg2_s3_w[1 ]), .i1(stg2_c3_w[0 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[0 ]), .s(stg3_s2[1  ]), .c(stg3_c2[1  ]), .co(stg3_co2[1  ]));
counter_5to3 u_a32_2  (.i0(stg2_s3_w[2 ]), .i1(stg2_c3_w[1 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[1 ]), .s(stg3_s2[2  ]), .c(stg3_c2[2  ]), .co(stg3_co2[2  ]));
counter_5to3 u_a32_3  (.i0(stg2_s3_w[3 ]), .i1(stg2_c3_w[2 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[2 ]), .s(stg3_s2[3  ]), .c(stg3_c2[3  ]), .co(stg3_co2[3  ]));
counter_5to3 u_a32_4  (.i0(stg2_s3_w[4 ]), .i1(stg2_c3_w[3 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[3 ]), .s(stg3_s2[4  ]), .c(stg3_c2[4  ]), .co(stg3_co2[4  ]));
counter_5to3 u_a32_5  (.i0(stg2_s3_w[5 ]), .i1(stg2_c3_w[4 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[4 ]), .s(stg3_s2[5  ]), .c(stg3_c2[5  ]), .co(stg3_co2[5  ]));
counter_5to3 u_a32_6  (.i0(stg2_s3_w[6 ]), .i1(stg2_c3_w[5 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[5 ]), .s(stg3_s2[6  ]), .c(stg3_c2[6  ]), .co(stg3_co2[6  ]));
counter_5to3 u_a32_7  (.i0(stg2_s3_w[7 ]), .i1(stg2_c3_w[6 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[6 ]), .s(stg3_s2[7  ]), .c(stg3_c2[7  ]), .co(stg3_co2[7  ]));
counter_5to3 u_a32_8  (.i0(stg2_s3_w[8 ]), .i1(stg2_c3_w[7 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[7 ]), .s(stg3_s2[8  ]), .c(stg3_c2[8  ]), .co(stg3_co2[8  ]));
counter_5to3 u_a32_9  (.i0(stg2_s3_w[9 ]), .i1(stg2_c3_w[8 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[8 ]), .s(stg3_s2[9  ]), .c(stg3_c2[9  ]), .co(stg3_co2[9  ]));
counter_5to3 u_a32_10 (.i0(stg2_s3_w[10]), .i1(stg2_c3_w[9 ]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[9 ]), .s(stg3_s2[10 ]), .c(stg3_c2[10 ]), .co(stg3_co2[10 ]));
counter_5to3 u_a32_11 (.i0(stg2_s3_w[11]), .i1(stg2_c3_w[10]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[10]), .s(stg3_s2[11 ]), .c(stg3_c2[11 ]), .co(stg3_co2[11 ]));
counter_5to3 u_a32_12 (.i0(stg2_s3_w[12]), .i1(stg2_c3_w[11]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[11]), .s(stg3_s2[12 ]), .c(stg3_c2[12 ]), .co(stg3_co2[12 ]));
counter_5to3 u_a32_13 (.i0(stg2_s3_w[13]), .i1(stg2_c3_w[12]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[12]), .s(stg3_s2[13 ]), .c(stg3_c2[13 ]), .co(stg3_co2[13 ]));
counter_5to3 u_a32_14 (.i0(stg2_s3_w[14]), .i1(stg2_c3_w[13]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[13]), .s(stg3_s2[14 ]), .c(stg3_c2[14 ]), .co(stg3_co2[14 ]));
counter_5to3 u_a32_15 (.i0(stg2_s3_w[15]), .i1(stg2_c3_w[14]), .i2(1'b0         ), .i3(1'b0         ), .ci(stg3_co2[14]), .s(stg3_s2[15 ]), .c(stg3_c2[15 ]), .co(stg3_co2[15 ]));
counter_5to3 u_a32_16 (.i0(stg2_s3_w[16]), .i1(stg2_c3_w[15]), .i2(stg2_s4_w[0 ]), .i3(1'b0         ), .ci(stg3_co2[15]), .s(stg3_s2[16 ]), .c(stg3_c2[16 ]), .co(stg3_co2[16 ]));
counter_5to3 u_a32_17 (.i0(stg2_s3_w[17]), .i1(stg2_c3_w[16]), .i2(stg2_s4_w[1 ]), .i3(stg2_c4_w[0 ]), .ci(stg3_co2[16]), .s(stg3_s2[17 ]), .c(stg3_c2[17 ]), .co(stg3_co2[17 ]));
counter_5to3 u_a32_18 (.i0(stg2_s3_w[18]), .i1(stg2_c3_w[17]), .i2(stg2_s4_w[2 ]), .i3(stg2_c4_w[1 ]), .ci(stg3_co2[17]), .s(stg3_s2[18 ]), .c(stg3_c2[18 ]), .co(stg3_co2[18 ]));
counter_5to3 u_a32_19 (.i0(stg2_s3_w[19]), .i1(stg2_c3_w[18]), .i2(stg2_s4_w[3 ]), .i3(stg2_c4_w[2 ]), .ci(stg3_co2[18]), .s(stg3_s2[19 ]), .c(stg3_c2[19 ]), .co(stg3_co2[19 ]));
counter_5to3 u_a32_20 (.i0(stg2_s3_w[20]), .i1(stg2_c3_w[19]), .i2(stg2_s4_w[4 ]), .i3(stg2_c4_w[3 ]), .ci(stg3_co2[19]), .s(stg3_s2[20 ]), .c(stg3_c2[20 ]), .co(stg3_co2[20 ]));
counter_5to3 u_a32_21 (.i0(stg2_s3_w[21]), .i1(stg2_c3_w[20]), .i2(stg2_s4_w[5 ]), .i3(stg2_c4_w[4 ]), .ci(stg3_co2[20]), .s(stg3_s2[21 ]), .c(stg3_c2[21 ]), .co(stg3_co2[21 ]));
counter_5to3 u_a32_22 (.i0(stg2_s3_w[22]), .i1(stg2_c3_w[21]), .i2(stg2_s4_w[6 ]), .i3(stg2_c4_w[5 ]), .ci(stg3_co2[21]), .s(stg3_s2[22 ]), .c(stg3_c2[22 ]), .co(stg3_co2[22 ]));
counter_5to3 u_a32_23 (.i0(stg2_s3_w[23]), .i1(stg2_c3_w[22]), .i2(stg2_s4_w[7 ]), .i3(stg2_c4_w[6 ]), .ci(stg3_co2[22]), .s(stg3_s2[23 ]), .c(stg3_c2[23 ]), .co(stg3_co2[23 ]));
counter_5to3 u_a32_24 (.i0(stg2_s3_w[24]), .i1(stg2_c3_w[23]), .i2(stg2_s4_w[8 ]), .i3(stg2_c4_w[7 ]), .ci(stg3_co2[23]), .s(stg3_s2[24 ]), .c(stg3_c2[24 ]), .co(stg3_co2[24 ]));
counter_5to3 u_a32_25 (.i0(stg2_s3_w[25]), .i1(stg2_c3_w[24]), .i2(stg2_s4_w[9 ]), .i3(stg2_c4_w[8 ]), .ci(stg3_co2[24]), .s(stg3_s2[25 ]), .c(stg3_c2[25 ]), .co(stg3_co2[25 ]));
counter_5to3 u_a32_26 (.i0(stg2_s3_w[26]), .i1(stg2_c3_w[25]), .i2(stg2_s4_w[10]), .i3(stg2_c4_w[9 ]), .ci(stg3_co2[25]), .s(stg3_s2[26 ]), .c(stg3_c2[26 ]), .co(stg3_co2[26 ]));
counter_5to3 u_a32_27 (.i0(stg2_s3_w[27]), .i1(stg2_c3_w[26]), .i2(stg2_s4_w[11]), .i3(stg2_c4_w[10]), .ci(stg3_co2[26]), .s(stg3_s2[27 ]), .c(stg3_c2[27 ]), .co(stg3_co2[27 ]));
counter_5to3 u_a32_28 (.i0(stg2_s3_w[28]), .i1(stg2_c3_w[27]), .i2(stg2_s4_w[12]), .i3(stg2_c4_w[11]), .ci(stg3_co2[27]), .s(stg3_s2[28 ]), .c(stg3_c2[28 ]), .co(stg3_co2[28 ]));
counter_5to3 u_a32_29 (.i0(stg2_s3_w[29]), .i1(stg2_c3_w[28]), .i2(stg2_s4_w[13]), .i3(stg2_c4_w[12]), .ci(stg3_co2[28]), .s(stg3_s2[29 ]), .c(stg3_c2[29 ]), .co(stg3_co2[29 ]));
counter_5to3 u_a32_30 (.i0(stg2_s3_w[30]), .i1(stg2_c3_w[29]), .i2(stg2_s4_w[14]), .i3(stg2_c4_w[13]), .ci(stg3_co2[29]), .s(stg3_s2[30 ]), .c(stg3_c2[30 ]), .co(stg3_co2[30 ]));
counter_5to3 u_a32_31 (.i0(stg2_s3_w[31]), .i1(stg2_c3_w[30]), .i2(stg2_s4_w[15]), .i3(stg2_c4_w[14]), .ci(stg3_co2[30]), .s(stg3_s2[31 ]), .c(stg3_c2[31 ]), .co(stg3_co2[31 ]));
counter_5to3 u_a32_32 (.i0(stg2_s3_w[32]), .i1(stg2_c3_w[31]), .i2(stg2_s4_w[16]), .i3(stg2_c4_w[15]), .ci(stg3_co2[31]), .s(stg3_s2[32 ]), .c(stg3_c2[32 ]), .co(stg3_co2[32 ]));
counter_5to3 u_a32_33 (.i0(stg2_s3_w[33]), .i1(stg2_c3_w[32]), .i2(stg2_s4_w[17]), .i3(stg2_c4_w[16]), .ci(stg3_co2[32]), .s(stg3_s2[33 ]), .c(stg3_c2[33 ]), .co(stg3_co2[33 ]));
counter_5to3 u_a32_34 (.i0(stg2_s3_w[34]), .i1(stg2_c3_w[33]), .i2(stg2_s4_w[18]), .i3(stg2_c4_w[17]), .ci(stg3_co2[33]), .s(stg3_s2[34 ]), .c(stg3_c2[34 ]), .co(stg3_co2[34 ]));
counter_5to3 u_a32_35 (.i0(stg2_s3_w[35]), .i1(stg2_c3_w[34]), .i2(stg2_s4_w[19]), .i3(stg2_c4_w[18]), .ci(stg3_co2[34]), .s(stg3_s2[35 ]), .c(stg3_c2[35 ]), .co(stg3_co2[35 ]));
counter_5to3 u_a32_36 (.i0(stg2_s3_w[36]), .i1(stg2_c3_w[35]), .i2(stg2_s4_w[20]), .i3(stg2_c4_w[19]), .ci(stg3_co2[35]), .s(stg3_s2[36 ]), .c(stg3_c2[36 ]), .co(stg3_co2[36 ]));
counter_5to3 u_a32_37 (.i0(stg2_s3_w[37]), .i1(stg2_c3_w[36]), .i2(stg2_s4_w[21]), .i3(stg2_c4_w[20]), .ci(stg3_co2[36]), .s(stg3_s2[37 ]), .c(stg3_c2[37 ]), .co(stg3_co2[37 ]));
counter_5to3 u_a32_38 (.i0(stg2_s3_w[38]), .i1(stg2_c3_w[37]), .i2(stg2_s4_w[22]), .i3(stg2_c4_w[21]), .ci(stg3_co2[37]), .s(stg3_s2[38 ]), .c(stg3_c2[38 ]), .co(stg3_co2[38 ]));
counter_5to3 u_a32_39 (.i0(stg2_s3_w[39]), .i1(stg2_c3_w[38]), .i2(stg2_s4_w[23]), .i3(stg2_c4_w[22]), .ci(stg3_co2[38]), .s(stg3_s2[39 ]), .c(stg3_c2[39 ]), .co(stg3_co2[39 ]));
counter_5to3 u_a32_40 (.i0(stg2_s3_w[40]), .i1(stg2_c3_w[39]), .i2(stg2_s4_w[24]), .i3(stg2_c4_w[23]), .ci(stg3_co2[39]), .s(stg3_s2[40 ]), .c(stg3_c2[40 ]), .co(stg3_co2[40 ]));
counter_5to3 u_a32_41 (.i0(stg2_s3_w[41]), .i1(stg2_c3_w[40]), .i2(stg2_s4_w[25]), .i3(stg2_c4_w[24]), .ci(stg3_co2[40]), .s(stg3_s2[41 ]), .c(stg3_c2[41 ]), .co(stg3_co2[41 ]));
counter_5to3 u_a32_42 (.i0(stg2_s3_w[42]), .i1(stg2_c3_w[41]), .i2(stg2_s4_w[26]), .i3(stg2_c4_w[25]), .ci(stg3_co2[41]), .s(stg3_s2[42 ]), .c(stg3_c2[42 ]), .co(stg3_co2[42 ]));
counter_5to3 u_a32_43 (.i0(stg2_s3_w[43]), .i1(stg2_c3_w[42]), .i2(stg2_s4_w[27]), .i3(stg2_c4_w[26]), .ci(stg3_co2[42]), .s(stg3_s2[43 ]), .c(stg3_c2[43 ]), .co(stg3_co2[43 ]));
counter_5to3 u_a32_44 (.i0(stg2_s3_w[44]), .i1(stg2_c3_w[43]), .i2(stg2_s4_w[28]), .i3(stg2_c4_w[27]), .ci(stg3_co2[43]), .s(stg3_s2[44 ]), .c(stg3_c2[44 ]), .co(stg3_co2[44 ]));
counter_5to3 u_a32_45 (.i0(stg2_s3_w[45]), .i1(stg2_c3_w[44]), .i2(stg2_s4_w[29]), .i3(stg2_c4_w[28]), .ci(stg3_co2[44]), .s(stg3_s2[45 ]), .c(stg3_c2[45 ]), .co(stg3_co2[45 ]));
counter_5to3 u_a32_46 (.i0(stg2_s3_w[46]), .i1(stg2_c3_w[45]), .i2(stg2_s4_w[30]), .i3(stg2_c4_w[29]), .ci(stg3_co2[45]), .s(stg3_s2[46 ]), .c(stg3_c2[46 ]), .co(stg3_co2[46 ]));
counter_5to3 u_a32_47 (.i0(stg2_s3_w[47]), .i1(stg2_c3_w[46]), .i2(stg2_s4_w[31]), .i3(stg2_c4_w[30]), .ci(stg3_co2[46]), .s(stg3_s2[47 ]), .c(stg3_c2[47 ]), .co(stg3_co2[47 ]));
counter_5to3 u_a32_48 (.i0(stg2_s3_w[48]), .i1(stg2_c3_w[47]), .i2(stg2_s4_w[32]), .i3(stg2_c4_w[31]), .ci(stg3_co2[47]), .s(stg3_s2[48 ]), .c(stg3_c2[48 ]), .co(stg3_co2[48 ]));
counter_5to3 u_a32_49 (.i0(stg2_s3_w[49]), .i1(stg2_c3_w[48]), .i2(stg2_s4_w[33]), .i3(stg2_c4_w[32]), .ci(stg3_co2[48]), .s(stg3_s2[49 ]), .c(stg3_c2[49 ]), .co(stg3_co2[49 ]));
counter_5to3 u_a32_50 (.i0(stg2_s3_w[50]), .i1(stg2_c3_w[49]), .i2(stg2_s4_w[34]), .i3(stg2_c4_w[33]), .ci(stg3_co2[49]), .s(stg3_s2[50 ]), .c(stg3_c2[50 ]), .co(stg3_co2[50 ]));
counter_5to3 u_a32_51 (.i0(stg2_s3_w[51]), .i1(stg2_c3_w[50]), .i2(stg2_s4_w[35]), .i3(stg2_c4_w[34]), .ci(stg3_co2[50]), .s(stg3_s2[51 ]), .c(stg3_c2[51 ]), .co(stg3_co2[51 ]));
counter_5to3 u_a32_52 (.i0(stg2_s3_w[52]), .i1(stg2_c3_w[51]), .i2(stg2_s4_w[36]), .i3(stg2_c4_w[35]), .ci(stg3_co2[51]), .s(stg3_s2[52 ]), .c(stg3_c2[52 ]), .co(stg3_co2[52 ]));
counter_5to3 u_a32_53 (.i0(stg2_s3_w[53]), .i1(stg2_c3_w[52]), .i2(stg2_s4_w[37]), .i3(stg2_c4_w[36]), .ci(stg3_co2[52]), .s(stg3_s2[53 ]), .c(stg3_c2[53 ]), .co(stg3_co2[53 ]));
counter_5to3 u_a32_54 (.i0(stg2_s3_w[54]), .i1(stg2_c3_w[53]), .i2(stg2_s4_w[38]), .i3(stg2_c4_w[37]), .ci(stg3_co2[53]), .s(stg3_s2[54 ]), .c(stg3_c2[54 ]), .co(stg3_co2[54 ]));
counter_5to3 u_a32_55 (.i0(stg2_s3_w[55]), .i1(stg2_c3_w[54]), .i2(stg2_s4_w[39]), .i3(stg2_c4_w[38]), .ci(stg3_co2[54]), .s(stg3_s2[55 ]), .c(stg3_c2[55 ]), .co(stg3_co2[55 ]));
counter_5to3 u_a32_56 (.i0(stg2_s3_w[56]), .i1(stg2_c3_w[55]), .i2(stg2_s4_w[40]), .i3(stg2_c4_w[39]), .ci(stg3_co2[55]), .s(stg3_s2[56 ]), .c(stg3_c2[56 ]), .co(stg3_co2[56 ]));
counter_5to3 u_a32_57 (.i0(stg2_s3_w[57]), .i1(stg2_c3_w[56]), .i2(stg2_s4_w[41]), .i3(stg2_c4_w[40]), .ci(stg3_co2[56]), .s(stg3_s2[57 ]), .c(stg3_c2[57 ]), .co(stg3_co2[57 ]));
counter_5to3 u_a32_58 (.i0(stg2_s3_w[58]), .i1(stg2_c3_w[57]), .i2(stg2_s4_w[42]), .i3(stg2_c4_w[41]), .ci(stg3_co2[57]), .s(stg3_s2[58 ]), .c(stg3_c2[58 ]), .co(stg3_co2[58 ]));
counter_5to3 u_a32_59 (.i0(stg2_s3_w[59]), .i1(stg2_c3_w[58]), .i2(stg2_s4_w[43]), .i3(stg2_c4_w[42]), .ci(stg3_co2[58]), .s(stg3_s2[59 ]), .c(stg3_c2[59 ]), .co(stg3_co2[59 ]));
counter_5to3 u_a32_60 (.i0(stg2_s3_w[60]), .i1(stg2_c3_w[59]), .i2(stg2_s4_w[44]), .i3(stg2_c4_w[43]), .ci(stg3_co2[59]), .s(stg3_s2[60 ]), .c(stg3_c2[60 ]), .co(stg3_co2[60 ]));
counter_5to3 u_a32_61 (.i0(stg2_s3_w[61]), .i1(stg2_c3_w[60]), .i2(stg2_s4_w[45]), .i3(stg2_c4_w[44]), .ci(stg3_co2[60]), .s(stg3_s2[61 ]), .c(stg3_c2[61 ]), .co(stg3_co2[61 ]));
counter_5to3 u_a32_62 (.i0(stg2_s3_w[62]), .i1(stg2_c3_w[61]), .i2(stg2_s4_w[46]), .i3(stg2_c4_w[45]), .ci(stg3_co2[61]), .s(stg3_s2[62 ]), .c(stg3_c2[62 ]), .co(stg3_co2[62 ]));
counter_5to3 u_a32_63 (.i0(stg2_s3_w[63]), .i1(stg2_c3_w[62]), .i2(stg2_s4_w[47]), .i3(stg2_c4_w[46]), .ci(stg3_co2[62]), .s(stg3_s2[63 ]), .c(stg3_c2[63 ]), .co(stg3_co2[63 ]));
counter_5to3 u_a32_64 (.i0(stg2_s3_w[64]), .i1(stg2_c3_w[63]), .i2(stg2_s4_w[48]), .i3(stg2_c4_w[47]), .ci(stg3_co2[63]), .s(stg3_s2[64 ]), .c(stg3_c2[64 ]), .co(stg3_co2[64 ]));
counter_5to3 u_a32_65 (.i0(stg2_s3_w[65]), .i1(stg2_c3_w[64]), .i2(stg2_s4_w[49]), .i3(stg2_c4_w[48]), .ci(stg3_co2[64]), .s(stg3_s2[65 ]), .c(stg3_c2[65 ]), .co(stg3_co2[65 ]));
counter_5to3 u_a32_66 (.i0(stg2_s3_w[66]), .i1(stg2_c3_w[65]), .i2(stg2_s4_w[50]), .i3(stg2_c4_w[49]), .ci(stg3_co2[65]), .s(stg3_s2[66 ]), .c(stg3_c2[66 ]), .co(stg3_co2[66 ]));
counter_5to3 u_a32_67 (.i0(stg2_s3_w[67]), .i1(stg2_c3_w[66]), .i2(stg2_s4_w[51]), .i3(stg2_c4_w[50]), .ci(stg3_co2[66]), .s(stg3_s2[67 ]), .c(stg3_c2[67 ]), .co(stg3_co2[67 ]));
counter_5to3 u_a32_68 (.i0(stg2_s3_w[68]), .i1(stg2_c3_w[67]), .i2(stg2_s4_w[52]), .i3(stg2_c4_w[51]), .ci(stg3_co2[67]), .s(stg3_s2[68 ]), .c(stg3_c2[68 ]), .co(stg3_co2[68 ]));
counter_5to3 u_a32_69 (.i0(stg2_s3_w[69]), .i1(stg2_c3_w[68]), .i2(stg2_s4_w[53]), .i3(stg2_c4_w[52]), .ci(stg3_co2[68]), .s(stg3_s2[69 ]), .c(stg3_c2[69 ]), .co(stg3_co2[69 ]));
counter_5to3 u_a32_70 (.i0(stg2_s3_w[70]), .i1(stg2_c3_w[69]), .i2(stg2_s4_w[54]), .i3(stg2_c4_w[53]), .ci(stg3_co2[69]), .s(stg3_s2[70 ]), .c(stg3_c2[70 ]), .co(stg3_co2[70 ]));
counter_5to3 u_a32_71 (.i0(stg2_s3_w[71]), .i1(stg2_c3_w[70]), .i2(stg2_s4_w[55]), .i3(stg2_c4_w[54]), .ci(stg3_co2[70]), .s(stg3_s2[71 ]), .c(stg3_c2[71 ]), .co(stg3_co2[71 ]));
counter_5to3 u_a32_72 (.i0(stg2_s3_w[72]), .i1(stg2_c3_w[71]), .i2(stg2_s4_w[56]), .i3(stg2_c4_w[55]), .ci(stg3_co2[71]), .s(stg3_s2[72 ]), .c(stg3_c2[72 ]), .co(stg3_co2[72 ]));
counter_5to3 u_a32_73 (.i0(stg2_s3_w[73]), .i1(stg2_c3_w[72]), .i2(stg2_s4_w[57]), .i3(stg2_c4_w[56]), .ci(stg3_co2[72]), .s(stg3_s2[73 ]), .c(stg3_c2[73 ]), .co(stg3_co2[73 ]));
counter_5to3 u_a32_74 (.i0(stg2_s3_w[74]), .i1(stg2_c3_w[73]), .i2(stg2_s4_w[58]), .i3(stg2_c4_w[57]), .ci(stg3_co2[73]), .s(stg3_s2[74 ]), .c(stg3_c2[74 ]), .co(stg3_co2[74 ]));
counter_5to3 u_a32_75 (.i0(stg2_s3_w[75]), .i1(stg2_c3_w[74]), .i2(stg2_s4_w[59]), .i3(stg2_c4_w[58]), .ci(stg3_co2[74]), .s(stg3_s2[75 ]), .c(stg3_c2[75 ]), .co(stg3_co2[75 ]));
counter_5to3 u_a32_76 (.i0(stg2_s3_w[76]), .i1(stg2_c3_w[75]), .i2(stg2_s4_w[60]), .i3(stg2_c4_w[59]), .ci(stg3_co2[75]), .s(stg3_s2[76 ]), .c(stg3_c2[76 ]), .co(stg3_co2[76 ]));
counter_5to3 u_a32_77 (.i0(stg2_s3_w[77]), .i1(stg2_c3_w[76]), .i2(stg2_s4_w[61]), .i3(stg2_c4_w[60]), .ci(stg3_co2[76]), .s(stg3_s2[77 ]), .c(stg3_c2[77 ]), .co(stg3_co2[77 ]));
counter_5to3 u_a32_78 (.i0(stg2_s3_w[78]), .i1(stg2_c3_w[77]), .i2(stg2_s4_w[62]), .i3(stg2_c4_w[61]), .ci(stg3_co2[77]), .s(stg3_s2[78 ]), .c(stg3_c2[78 ]), .co(stg3_co2[78 ]));
counter_5to3 u_a32_79 (.i0(stg2_s3_w[79]), .i1(stg2_c3_w[78]), .i2(stg2_s4_w[63]), .i3(stg2_c4_w[62]), .ci(stg3_co2[78]), .s(stg3_s2[79 ]), .c(stg3_c2[79 ]), .co(stg3_co2[79 ]));
counter_5to3 u_a32_80 (.i0(stg2_s3_w[80]), .i1(stg2_c3_w[79]), .i2(stg2_s4_w[64]), .i3(stg2_c4_w[63]), .ci(stg3_co2[79]), .s(stg3_s2[80 ]), .c(stg3_c2[80 ]), .co(stg3_co2[80 ]));
counter_5to3 u_a32_81 (.i0(stg2_s3_w[81]), .i1(stg2_c3_w[80]), .i2(stg2_s4_w[65]), .i3(stg2_c4_w[64]), .ci(stg3_co2[80]), .s(stg3_s2[81 ]), .c(stg3_c2[81 ]), .co(stg3_co2[81 ]));
counter_5to3 u_a32_82 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[81]), .i2(stg2_s4_w[66]), .i3(stg2_c4_w[65]), .ci(stg3_co2[81]), .s(stg3_s2[82 ]), .c(stg3_c2[82 ]), .co(stg3_co2[82 ]));
counter_5to3 u_a32_83 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[67]), .i3(stg2_c4_w[66]), .ci(stg3_co2[82]), .s(stg3_s2[83 ]), .c(stg3_c2[83 ]), .co(stg3_co2[83 ]));
counter_5to3 u_a32_84 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[68]), .i3(stg2_c4_w[67]), .ci(stg3_co2[83]), .s(stg3_s2[84 ]), .c(stg3_c2[84 ]), .co(stg3_co2[84 ]));
counter_5to3 u_a32_85 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[69]), .i3(stg2_c4_w[68]), .ci(stg3_co2[84]), .s(stg3_s2[85 ]), .c(stg3_c2[85 ]), .co(stg3_co2[85 ]));
counter_5to3 u_a32_86 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[70]), .i3(stg2_c4_w[69]), .ci(stg3_co2[85]), .s(stg3_s2[86 ]), .c(stg3_c2[86 ]), .co(stg3_co2[86 ]));
counter_5to3 u_a32_87 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[71]), .i3(stg2_c4_w[70]), .ci(stg3_co2[86]), .s(stg3_s2[87 ]), .c(stg3_c2[87 ]), .co(stg3_co2[87 ]));
counter_5to3 u_a32_88 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[72]), .i3(stg2_c4_w[71]), .ci(stg3_co2[87]), .s(stg3_s2[88 ]), .c(stg3_c2[88 ]), .co(stg3_co2[88 ]));
counter_5to3 u_a32_89 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[73]), .i3(stg2_c4_w[72]), .ci(stg3_co2[88]), .s(stg3_s2[89 ]), .c(stg3_c2[89 ]), .co(stg3_co2[89 ]));
counter_5to3 u_a32_90 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[74]), .i3(stg2_c4_w[73]), .ci(stg3_co2[89]), .s(stg3_s2[90 ]), .c(stg3_c2[90 ]), .co(stg3_co2[90 ]));
counter_5to3 u_a32_91 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[75]), .i3(stg2_c4_w[74]), .ci(stg3_co2[90]), .s(stg3_s2[91 ]), .c(stg3_c2[91 ]), .co(stg3_co2[91 ]));
counter_5to3 u_a32_92 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[76]), .i3(stg2_c4_w[75]), .ci(stg3_co2[91]), .s(stg3_s2[92 ]), .c(stg3_c2[92 ]), .co(stg3_co2[92 ]));
counter_5to3 u_a32_93 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[77]), .i3(stg2_c4_w[76]), .ci(stg3_co2[92]), .s(stg3_s2[93 ]), .c(stg3_c2[93 ]), .co(stg3_co2[93 ]));
counter_5to3 u_a32_94 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[78]), .i3(stg2_c4_w[77]), .ci(stg3_co2[93]), .s(stg3_s2[94 ]), .c(stg3_c2[94 ]), .co(stg3_co2[94 ]));
counter_5to3 u_a32_95 (.i0(stg2_s3_w[82]), .i1(stg2_c3_w[82]), .i2(stg2_s4_w[79]), .i3(stg2_c4_w[78]), .ci(stg3_co2[94]), .s(stg3_s2[95 ]), .c(stg3_c2[95 ]), .co(stg3_co2[95 ]));

//================ forth stage ================
wire [100:0] stg3_s1_w, stg3_c1_w;
wire [95:0] stg3_s2_w, stg3_c2_w;
wire [65:0] pp33_w3;

// ========= pipeline ============
reg [100:0] stg3_s1_ff, stg3_c1_ff;
reg [95:0]  stg3_s2_ff, stg3_c2_ff;
reg [65:0]  pp33_f3;

always @(posedge clk or negedge rstn)begin
    if (!rstn)begin
        stg3_s1_ff <= 101'b0;
        stg3_c1_ff <= 101'b0;
        stg3_s2_ff <= 96'b0;
        stg3_c2_ff <= 96'b0;
        pp33_f3    <= 66'b0;
    end
    else begin
        stg3_s1_ff <= stg3_s1;
        stg3_c1_ff <= stg3_c1;
        stg3_s2_ff <= stg3_s2;
        stg3_c2_ff <= stg3_c2;
        pp33_f3    <= pp33_w2;
    end
end

assign stg3_s1_w = stg3_s1_ff;
assign stg3_c1_w = stg3_c1_ff;
assign stg3_s2_w = stg3_s2_ff;
assign stg3_c2_w = stg3_c2_ff;
assign pp33_w3   = pp33_f3   ;


wire [127:0] stg4_s1, stg4_c1, stg4_co1;

// =========================== forth stage 1st group ============================================================================================================
counter_5to3 u_a41_0  (.i0(stg3_s1_w[0  ]), .i1(1'b0         ), .i2(1'b0         ), .i3(1'b0            ), .ci(1'b0         ), .s(stg4_s1[0  ]), .c(stg4_c1[0  ]), .co(stg4_co1[0  ]));
counter_5to3 u_a41_1  (.i0(stg3_s1_w[1  ]), .i1(stg3_c1_w[0  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[0  ]), .s(stg4_s1[1  ]), .c(stg4_c1[1  ]), .co(stg4_co1[1  ]));
counter_5to3 u_a41_2  (.i0(stg3_s1_w[2  ]), .i1(stg3_c1_w[1  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[1  ]), .s(stg4_s1[2  ]), .c(stg4_c1[2  ]), .co(stg4_co1[2  ]));
counter_5to3 u_a41_3  (.i0(stg3_s1_w[3  ]), .i1(stg3_c1_w[2  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[2  ]), .s(stg4_s1[3  ]), .c(stg4_c1[3  ]), .co(stg4_co1[3  ]));
counter_5to3 u_a41_4  (.i0(stg3_s1_w[4  ]), .i1(stg3_c1_w[3  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[3  ]), .s(stg4_s1[4  ]), .c(stg4_c1[4  ]), .co(stg4_co1[4  ]));
counter_5to3 u_a41_5  (.i0(stg3_s1_w[5  ]), .i1(stg3_c1_w[4  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[4  ]), .s(stg4_s1[5  ]), .c(stg4_c1[5  ]), .co(stg4_co1[5  ]));
counter_5to3 u_a41_6  (.i0(stg3_s1_w[6  ]), .i1(stg3_c1_w[5  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[5  ]), .s(stg4_s1[6  ]), .c(stg4_c1[6  ]), .co(stg4_co1[6  ]));
counter_5to3 u_a41_7  (.i0(stg3_s1_w[7  ]), .i1(stg3_c1_w[6  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[6  ]), .s(stg4_s1[7  ]), .c(stg4_c1[7  ]), .co(stg4_co1[7  ]));
counter_5to3 u_a41_8  (.i0(stg3_s1_w[8  ]), .i1(stg3_c1_w[7  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[7  ]), .s(stg4_s1[8  ]), .c(stg4_c1[8  ]), .co(stg4_co1[8  ]));
counter_5to3 u_a41_9  (.i0(stg3_s1_w[9  ]), .i1(stg3_c1_w[8  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[8  ]), .s(stg4_s1[9  ]), .c(stg4_c1[9  ]), .co(stg4_co1[9  ]));
counter_5to3 u_a41_10 (.i0(stg3_s1_w[10 ]), .i1(stg3_c1_w[9  ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[9  ]), .s(stg4_s1[10 ]), .c(stg4_c1[10 ]), .co(stg4_co1[10 ]));
counter_5to3 u_a41_11 (.i0(stg3_s1_w[11 ]), .i1(stg3_c1_w[10 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[10 ]), .s(stg4_s1[11 ]), .c(stg4_c1[11 ]), .co(stg4_co1[11 ]));
counter_5to3 u_a41_12 (.i0(stg3_s1_w[12 ]), .i1(stg3_c1_w[11 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[11 ]), .s(stg4_s1[12 ]), .c(stg4_c1[12 ]), .co(stg4_co1[12 ]));
counter_5to3 u_a41_13 (.i0(stg3_s1_w[13 ]), .i1(stg3_c1_w[12 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[12 ]), .s(stg4_s1[13 ]), .c(stg4_c1[13 ]), .co(stg4_co1[13 ]));
counter_5to3 u_a41_14 (.i0(stg3_s1_w[14 ]), .i1(stg3_c1_w[13 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[13 ]), .s(stg4_s1[14 ]), .c(stg4_c1[14 ]), .co(stg4_co1[14 ]));
counter_5to3 u_a41_15 (.i0(stg3_s1_w[15 ]), .i1(stg3_c1_w[14 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[14 ]), .s(stg4_s1[15 ]), .c(stg4_c1[15 ]), .co(stg4_co1[15 ]));
counter_5to3 u_a41_16 (.i0(stg3_s1_w[16 ]), .i1(stg3_c1_w[15 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[15 ]), .s(stg4_s1[16 ]), .c(stg4_c1[16 ]), .co(stg4_co1[16 ]));
counter_5to3 u_a41_17 (.i0(stg3_s1_w[17 ]), .i1(stg3_c1_w[16 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[16 ]), .s(stg4_s1[17 ]), .c(stg4_c1[17 ]), .co(stg4_co1[17 ]));
counter_5to3 u_a41_18 (.i0(stg3_s1_w[18 ]), .i1(stg3_c1_w[17 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[17 ]), .s(stg4_s1[18 ]), .c(stg4_c1[18 ]), .co(stg4_co1[18 ]));
counter_5to3 u_a41_19 (.i0(stg3_s1_w[19 ]), .i1(stg3_c1_w[18 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[18 ]), .s(stg4_s1[19 ]), .c(stg4_c1[19 ]), .co(stg4_co1[19 ]));
counter_5to3 u_a41_20 (.i0(stg3_s1_w[20 ]), .i1(stg3_c1_w[19 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[19 ]), .s(stg4_s1[20 ]), .c(stg4_c1[20 ]), .co(stg4_co1[20 ]));
counter_5to3 u_a41_21 (.i0(stg3_s1_w[21 ]), .i1(stg3_c1_w[20 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[20 ]), .s(stg4_s1[21 ]), .c(stg4_c1[21 ]), .co(stg4_co1[21 ]));
counter_5to3 u_a41_22 (.i0(stg3_s1_w[22 ]), .i1(stg3_c1_w[21 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[21 ]), .s(stg4_s1[22 ]), .c(stg4_c1[22 ]), .co(stg4_co1[22 ]));
counter_5to3 u_a41_23 (.i0(stg3_s1_w[23 ]), .i1(stg3_c1_w[22 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[22 ]), .s(stg4_s1[23 ]), .c(stg4_c1[23 ]), .co(stg4_co1[23 ]));
counter_5to3 u_a41_24 (.i0(stg3_s1_w[24 ]), .i1(stg3_c1_w[23 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[23 ]), .s(stg4_s1[24 ]), .c(stg4_c1[24 ]), .co(stg4_co1[24 ]));
counter_5to3 u_a41_25 (.i0(stg3_s1_w[25 ]), .i1(stg3_c1_w[24 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[24 ]), .s(stg4_s1[25 ]), .c(stg4_c1[25 ]), .co(stg4_co1[25 ]));
counter_5to3 u_a41_26 (.i0(stg3_s1_w[26 ]), .i1(stg3_c1_w[25 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[25 ]), .s(stg4_s1[26 ]), .c(stg4_c1[26 ]), .co(stg4_co1[26 ]));
counter_5to3 u_a41_27 (.i0(stg3_s1_w[27 ]), .i1(stg3_c1_w[26 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[26 ]), .s(stg4_s1[27 ]), .c(stg4_c1[27 ]), .co(stg4_co1[27 ]));
counter_5to3 u_a41_28 (.i0(stg3_s1_w[28 ]), .i1(stg3_c1_w[27 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[27 ]), .s(stg4_s1[28 ]), .c(stg4_c1[28 ]), .co(stg4_co1[28 ]));
counter_5to3 u_a41_29 (.i0(stg3_s1_w[29 ]), .i1(stg3_c1_w[28 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[28 ]), .s(stg4_s1[29 ]), .c(stg4_c1[29 ]), .co(stg4_co1[29 ]));
counter_5to3 u_a41_30 (.i0(stg3_s1_w[30 ]), .i1(stg3_c1_w[29 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[29 ]), .s(stg4_s1[30 ]), .c(stg4_c1[30 ]), .co(stg4_co1[30 ]));
counter_5to3 u_a41_31 (.i0(stg3_s1_w[31 ]), .i1(stg3_c1_w[30 ]), .i2(1'b0         ), .i3(1'b0           ), .ci(stg4_co1[30 ]), .s(stg4_s1[31 ]), .c(stg4_c1[31 ]), .co(stg4_co1[31 ]));
counter_5to3 u_a41_32 (.i0(stg3_s1_w[32 ]), .i1(stg3_c1_w[31 ]), .i2(stg3_s2_w[0  ]), .i3(1'b0          ), .ci(stg4_co1[31 ]), .s(stg4_s1[32 ]), .c(stg4_c1[32 ]), .co(stg4_co1[32 ]));
counter_5to3 u_a41_33 (.i0(stg3_s1_w[33 ]), .i1(stg3_c1_w[32 ]), .i2(stg3_s2_w[1  ]), .i3(stg3_c2_w[0  ]), .ci(stg4_co1[32 ]), .s(stg4_s1[33 ]), .c(stg4_c1[33 ]), .co(stg4_co1[33 ]));
counter_5to3 u_a41_34 (.i0(stg3_s1_w[34 ]), .i1(stg3_c1_w[33 ]), .i2(stg3_s2_w[2  ]), .i3(stg3_c2_w[1  ]), .ci(stg4_co1[33 ]), .s(stg4_s1[34 ]), .c(stg4_c1[34 ]), .co(stg4_co1[34 ]));
counter_5to3 u_a41_35 (.i0(stg3_s1_w[35 ]), .i1(stg3_c1_w[34 ]), .i2(stg3_s2_w[3  ]), .i3(stg3_c2_w[2  ]), .ci(stg4_co1[34 ]), .s(stg4_s1[35 ]), .c(stg4_c1[35 ]), .co(stg4_co1[35 ]));
counter_5to3 u_a41_36 (.i0(stg3_s1_w[36 ]), .i1(stg3_c1_w[35 ]), .i2(stg3_s2_w[4  ]), .i3(stg3_c2_w[3  ]), .ci(stg4_co1[35 ]), .s(stg4_s1[36 ]), .c(stg4_c1[36 ]), .co(stg4_co1[36 ]));
counter_5to3 u_a41_37 (.i0(stg3_s1_w[37 ]), .i1(stg3_c1_w[36 ]), .i2(stg3_s2_w[5  ]), .i3(stg3_c2_w[4  ]), .ci(stg4_co1[36 ]), .s(stg4_s1[37 ]), .c(stg4_c1[37 ]), .co(stg4_co1[37 ]));
counter_5to3 u_a41_38 (.i0(stg3_s1_w[38 ]), .i1(stg3_c1_w[37 ]), .i2(stg3_s2_w[6  ]), .i3(stg3_c2_w[5  ]), .ci(stg4_co1[37 ]), .s(stg4_s1[38 ]), .c(stg4_c1[38 ]), .co(stg4_co1[38 ]));
counter_5to3 u_a41_39 (.i0(stg3_s1_w[39 ]), .i1(stg3_c1_w[38 ]), .i2(stg3_s2_w[7  ]), .i3(stg3_c2_w[6  ]), .ci(stg4_co1[38 ]), .s(stg4_s1[39 ]), .c(stg4_c1[39 ]), .co(stg4_co1[39 ]));
counter_5to3 u_a41_40 (.i0(stg3_s1_w[40 ]), .i1(stg3_c1_w[39 ]), .i2(stg3_s2_w[8  ]), .i3(stg3_c2_w[7  ]), .ci(stg4_co1[39 ]), .s(stg4_s1[40 ]), .c(stg4_c1[40 ]), .co(stg4_co1[40 ]));
counter_5to3 u_a41_41 (.i0(stg3_s1_w[41 ]), .i1(stg3_c1_w[40 ]), .i2(stg3_s2_w[9  ]), .i3(stg3_c2_w[8  ]), .ci(stg4_co1[40 ]), .s(stg4_s1[41 ]), .c(stg4_c1[41 ]), .co(stg4_co1[41 ]));
counter_5to3 u_a41_42 (.i0(stg3_s1_w[42 ]), .i1(stg3_c1_w[41 ]), .i2(stg3_s2_w[10 ]), .i3(stg3_c2_w[9  ]), .ci(stg4_co1[41 ]), .s(stg4_s1[42 ]), .c(stg4_c1[42 ]), .co(stg4_co1[42 ]));
counter_5to3 u_a41_43 (.i0(stg3_s1_w[43 ]), .i1(stg3_c1_w[42 ]), .i2(stg3_s2_w[11 ]), .i3(stg3_c2_w[10 ]), .ci(stg4_co1[42 ]), .s(stg4_s1[43 ]), .c(stg4_c1[43 ]), .co(stg4_co1[43 ]));
counter_5to3 u_a41_44 (.i0(stg3_s1_w[44 ]), .i1(stg3_c1_w[43 ]), .i2(stg3_s2_w[12 ]), .i3(stg3_c2_w[11 ]), .ci(stg4_co1[43 ]), .s(stg4_s1[44 ]), .c(stg4_c1[44 ]), .co(stg4_co1[44 ]));
counter_5to3 u_a41_45 (.i0(stg3_s1_w[45 ]), .i1(stg3_c1_w[44 ]), .i2(stg3_s2_w[13 ]), .i3(stg3_c2_w[12 ]), .ci(stg4_co1[44 ]), .s(stg4_s1[45 ]), .c(stg4_c1[45 ]), .co(stg4_co1[45 ]));
counter_5to3 u_a41_46 (.i0(stg3_s1_w[46 ]), .i1(stg3_c1_w[45 ]), .i2(stg3_s2_w[14 ]), .i3(stg3_c2_w[13 ]), .ci(stg4_co1[45 ]), .s(stg4_s1[46 ]), .c(stg4_c1[46 ]), .co(stg4_co1[46 ]));
counter_5to3 u_a41_47 (.i0(stg3_s1_w[47 ]), .i1(stg3_c1_w[46 ]), .i2(stg3_s2_w[15 ]), .i3(stg3_c2_w[14 ]), .ci(stg4_co1[46 ]), .s(stg4_s1[47 ]), .c(stg4_c1[47 ]), .co(stg4_co1[47 ]));
counter_5to3 u_a41_48 (.i0(stg3_s1_w[48 ]), .i1(stg3_c1_w[47 ]), .i2(stg3_s2_w[16 ]), .i3(stg3_c2_w[15 ]), .ci(stg4_co1[47 ]), .s(stg4_s1[48 ]), .c(stg4_c1[48 ]), .co(stg4_co1[48 ]));
counter_5to3 u_a41_49 (.i0(stg3_s1_w[49 ]), .i1(stg3_c1_w[48 ]), .i2(stg3_s2_w[17 ]), .i3(stg3_c2_w[16 ]), .ci(stg4_co1[48 ]), .s(stg4_s1[49 ]), .c(stg4_c1[49 ]), .co(stg4_co1[49 ]));
counter_5to3 u_a41_50 (.i0(stg3_s1_w[50 ]), .i1(stg3_c1_w[49 ]), .i2(stg3_s2_w[18 ]), .i3(stg3_c2_w[17 ]), .ci(stg4_co1[49 ]), .s(stg4_s1[50 ]), .c(stg4_c1[50 ]), .co(stg4_co1[50 ]));
counter_5to3 u_a41_51 (.i0(stg3_s1_w[51 ]), .i1(stg3_c1_w[50 ]), .i2(stg3_s2_w[19 ]), .i3(stg3_c2_w[18 ]), .ci(stg4_co1[50 ]), .s(stg4_s1[51 ]), .c(stg4_c1[51 ]), .co(stg4_co1[51 ]));
counter_5to3 u_a41_52 (.i0(stg3_s1_w[52 ]), .i1(stg3_c1_w[51 ]), .i2(stg3_s2_w[20 ]), .i3(stg3_c2_w[19 ]), .ci(stg4_co1[51 ]), .s(stg4_s1[52 ]), .c(stg4_c1[52 ]), .co(stg4_co1[52 ]));
counter_5to3 u_a41_53 (.i0(stg3_s1_w[53 ]), .i1(stg3_c1_w[52 ]), .i2(stg3_s2_w[21 ]), .i3(stg3_c2_w[20 ]), .ci(stg4_co1[52 ]), .s(stg4_s1[53 ]), .c(stg4_c1[53 ]), .co(stg4_co1[53 ]));
counter_5to3 u_a41_54 (.i0(stg3_s1_w[54 ]), .i1(stg3_c1_w[53 ]), .i2(stg3_s2_w[22 ]), .i3(stg3_c2_w[21 ]), .ci(stg4_co1[53 ]), .s(stg4_s1[54 ]), .c(stg4_c1[54 ]), .co(stg4_co1[54 ]));
counter_5to3 u_a41_55 (.i0(stg3_s1_w[55 ]), .i1(stg3_c1_w[54 ]), .i2(stg3_s2_w[23 ]), .i3(stg3_c2_w[22 ]), .ci(stg4_co1[54 ]), .s(stg4_s1[55 ]), .c(stg4_c1[55 ]), .co(stg4_co1[55 ]));
counter_5to3 u_a41_56 (.i0(stg3_s1_w[56 ]), .i1(stg3_c1_w[55 ]), .i2(stg3_s2_w[24 ]), .i3(stg3_c2_w[23 ]), .ci(stg4_co1[55 ]), .s(stg4_s1[56 ]), .c(stg4_c1[56 ]), .co(stg4_co1[56 ]));
counter_5to3 u_a41_57 (.i0(stg3_s1_w[57 ]), .i1(stg3_c1_w[56 ]), .i2(stg3_s2_w[25 ]), .i3(stg3_c2_w[24 ]), .ci(stg4_co1[56 ]), .s(stg4_s1[57 ]), .c(stg4_c1[57 ]), .co(stg4_co1[57 ]));
counter_5to3 u_a41_58 (.i0(stg3_s1_w[58 ]), .i1(stg3_c1_w[57 ]), .i2(stg3_s2_w[26 ]), .i3(stg3_c2_w[25 ]), .ci(stg4_co1[57 ]), .s(stg4_s1[58 ]), .c(stg4_c1[58 ]), .co(stg4_co1[58 ]));
counter_5to3 u_a41_59 (.i0(stg3_s1_w[59 ]), .i1(stg3_c1_w[58 ]), .i2(stg3_s2_w[27 ]), .i3(stg3_c2_w[26 ]), .ci(stg4_co1[58 ]), .s(stg4_s1[59 ]), .c(stg4_c1[59 ]), .co(stg4_co1[59 ]));
counter_5to3 u_a41_60 (.i0(stg3_s1_w[60 ]), .i1(stg3_c1_w[59 ]), .i2(stg3_s2_w[28 ]), .i3(stg3_c2_w[27 ]), .ci(stg4_co1[59 ]), .s(stg4_s1[60 ]), .c(stg4_c1[60 ]), .co(stg4_co1[60 ]));
counter_5to3 u_a41_61 (.i0(stg3_s1_w[61 ]), .i1(stg3_c1_w[60 ]), .i2(stg3_s2_w[29 ]), .i3(stg3_c2_w[28 ]), .ci(stg4_co1[60 ]), .s(stg4_s1[61 ]), .c(stg4_c1[61 ]), .co(stg4_co1[61 ]));
counter_5to3 u_a41_62 (.i0(stg3_s1_w[62 ]), .i1(stg3_c1_w[61 ]), .i2(stg3_s2_w[30 ]), .i3(stg3_c2_w[29 ]), .ci(stg4_co1[61 ]), .s(stg4_s1[62 ]), .c(stg4_c1[62 ]), .co(stg4_co1[62 ]));
counter_5to3 u_a41_63 (.i0(stg3_s1_w[63 ]), .i1(stg3_c1_w[62 ]), .i2(stg3_s2_w[31 ]), .i3(stg3_c2_w[30 ]), .ci(stg4_co1[62 ]), .s(stg4_s1[63 ]), .c(stg4_c1[63 ]), .co(stg4_co1[63 ]));
counter_5to3 u_a41_64 (.i0(stg3_s1_w[64 ]), .i1(stg3_c1_w[63 ]), .i2(stg3_s2_w[32 ]), .i3(stg3_c2_w[31 ]), .ci(stg4_co1[63 ]), .s(stg4_s1[64 ]), .c(stg4_c1[64 ]), .co(stg4_co1[64 ]));
counter_5to3 u_a41_65 (.i0(stg3_s1_w[65 ]), .i1(stg3_c1_w[64 ]), .i2(stg3_s2_w[33 ]), .i3(stg3_c2_w[32 ]), .ci(stg4_co1[64 ]), .s(stg4_s1[65 ]), .c(stg4_c1[65 ]), .co(stg4_co1[65 ]));
counter_5to3 u_a41_66 (.i0(stg3_s1_w[66 ]), .i1(stg3_c1_w[65 ]), .i2(stg3_s2_w[34 ]), .i3(stg3_c2_w[33 ]), .ci(stg4_co1[65 ]), .s(stg4_s1[66 ]), .c(stg4_c1[66 ]), .co(stg4_co1[66 ]));
counter_5to3 u_a41_67 (.i0(stg3_s1_w[67 ]), .i1(stg3_c1_w[66 ]), .i2(stg3_s2_w[35 ]), .i3(stg3_c2_w[34 ]), .ci(stg4_co1[66 ]), .s(stg4_s1[67 ]), .c(stg4_c1[67 ]), .co(stg4_co1[67 ]));
counter_5to3 u_a41_68 (.i0(stg3_s1_w[68 ]), .i1(stg3_c1_w[67 ]), .i2(stg3_s2_w[36 ]), .i3(stg3_c2_w[35 ]), .ci(stg4_co1[67 ]), .s(stg4_s1[68 ]), .c(stg4_c1[68 ]), .co(stg4_co1[68 ]));
counter_5to3 u_a41_69 (.i0(stg3_s1_w[69 ]), .i1(stg3_c1_w[68 ]), .i2(stg3_s2_w[37 ]), .i3(stg3_c2_w[36 ]), .ci(stg4_co1[68 ]), .s(stg4_s1[69 ]), .c(stg4_c1[69 ]), .co(stg4_co1[69 ]));
counter_5to3 u_a41_70 (.i0(stg3_s1_w[70 ]), .i1(stg3_c1_w[69 ]), .i2(stg3_s2_w[38 ]), .i3(stg3_c2_w[37 ]), .ci(stg4_co1[69 ]), .s(stg4_s1[70 ]), .c(stg4_c1[70 ]), .co(stg4_co1[70 ]));
counter_5to3 u_a41_71 (.i0(stg3_s1_w[71 ]), .i1(stg3_c1_w[70 ]), .i2(stg3_s2_w[39 ]), .i3(stg3_c2_w[38 ]), .ci(stg4_co1[70 ]), .s(stg4_s1[71 ]), .c(stg4_c1[71 ]), .co(stg4_co1[71 ]));
counter_5to3 u_a41_72 (.i0(stg3_s1_w[72 ]), .i1(stg3_c1_w[71 ]), .i2(stg3_s2_w[40 ]), .i3(stg3_c2_w[39 ]), .ci(stg4_co1[71 ]), .s(stg4_s1[72 ]), .c(stg4_c1[72 ]), .co(stg4_co1[72 ]));
counter_5to3 u_a41_73 (.i0(stg3_s1_w[73 ]), .i1(stg3_c1_w[72 ]), .i2(stg3_s2_w[41 ]), .i3(stg3_c2_w[40 ]), .ci(stg4_co1[72 ]), .s(stg4_s1[73 ]), .c(stg4_c1[73 ]), .co(stg4_co1[73 ]));
counter_5to3 u_a41_74 (.i0(stg3_s1_w[74 ]), .i1(stg3_c1_w[73 ]), .i2(stg3_s2_w[42 ]), .i3(stg3_c2_w[41 ]), .ci(stg4_co1[73 ]), .s(stg4_s1[74 ]), .c(stg4_c1[74 ]), .co(stg4_co1[74 ]));
counter_5to3 u_a41_75 (.i0(stg3_s1_w[75 ]), .i1(stg3_c1_w[74 ]), .i2(stg3_s2_w[43 ]), .i3(stg3_c2_w[42 ]), .ci(stg4_co1[74 ]), .s(stg4_s1[75 ]), .c(stg4_c1[75 ]), .co(stg4_co1[75 ]));
counter_5to3 u_a41_76 (.i0(stg3_s1_w[76 ]), .i1(stg3_c1_w[75 ]), .i2(stg3_s2_w[44 ]), .i3(stg3_c2_w[43 ]), .ci(stg4_co1[75 ]), .s(stg4_s1[76 ]), .c(stg4_c1[76 ]), .co(stg4_co1[76 ]));
counter_5to3 u_a41_77 (.i0(stg3_s1_w[77 ]), .i1(stg3_c1_w[76 ]), .i2(stg3_s2_w[45 ]), .i3(stg3_c2_w[44 ]), .ci(stg4_co1[76 ]), .s(stg4_s1[77 ]), .c(stg4_c1[77 ]), .co(stg4_co1[77 ]));
counter_5to3 u_a41_78 (.i0(stg3_s1_w[78 ]), .i1(stg3_c1_w[77 ]), .i2(stg3_s2_w[46 ]), .i3(stg3_c2_w[45 ]), .ci(stg4_co1[77 ]), .s(stg4_s1[78 ]), .c(stg4_c1[78 ]), .co(stg4_co1[78 ]));
counter_5to3 u_a41_79 (.i0(stg3_s1_w[79 ]), .i1(stg3_c1_w[78 ]), .i2(stg3_s2_w[47 ]), .i3(stg3_c2_w[46 ]), .ci(stg4_co1[78 ]), .s(stg4_s1[79 ]), .c(stg4_c1[79 ]), .co(stg4_co1[79 ]));
counter_5to3 u_a41_80 (.i0(stg3_s1_w[80 ]), .i1(stg3_c1_w[79 ]), .i2(stg3_s2_w[48 ]), .i3(stg3_c2_w[47 ]), .ci(stg4_co1[79 ]), .s(stg4_s1[80 ]), .c(stg4_c1[80 ]), .co(stg4_co1[80 ]));
counter_5to3 u_a41_81 (.i0(stg3_s1_w[81 ]), .i1(stg3_c1_w[80 ]), .i2(stg3_s2_w[49 ]), .i3(stg3_c2_w[48 ]), .ci(stg4_co1[80 ]), .s(stg4_s1[81 ]), .c(stg4_c1[81 ]), .co(stg4_co1[81 ]));
counter_5to3 u_a41_82 (.i0(stg3_s1_w[82 ]), .i1(stg3_c1_w[81 ]), .i2(stg3_s2_w[50 ]), .i3(stg3_c2_w[49 ]), .ci(stg4_co1[81 ]), .s(stg4_s1[82 ]), .c(stg4_c1[82 ]), .co(stg4_co1[82 ]));
counter_5to3 u_a41_83 (.i0(stg3_s1_w[83 ]), .i1(stg3_c1_w[82 ]), .i2(stg3_s2_w[51 ]), .i3(stg3_c2_w[50 ]), .ci(stg4_co1[82 ]), .s(stg4_s1[83 ]), .c(stg4_c1[83 ]), .co(stg4_co1[83 ]));
counter_5to3 u_a41_84 (.i0(stg3_s1_w[84 ]), .i1(stg3_c1_w[83 ]), .i2(stg3_s2_w[52 ]), .i3(stg3_c2_w[51 ]), .ci(stg4_co1[83 ]), .s(stg4_s1[84 ]), .c(stg4_c1[84 ]), .co(stg4_co1[84 ]));
counter_5to3 u_a41_85 (.i0(stg3_s1_w[85 ]), .i1(stg3_c1_w[84 ]), .i2(stg3_s2_w[53 ]), .i3(stg3_c2_w[52 ]), .ci(stg4_co1[84 ]), .s(stg4_s1[85 ]), .c(stg4_c1[85 ]), .co(stg4_co1[85 ]));
counter_5to3 u_a41_86 (.i0(stg3_s1_w[86 ]), .i1(stg3_c1_w[85 ]), .i2(stg3_s2_w[54 ]), .i3(stg3_c2_w[53 ]), .ci(stg4_co1[85 ]), .s(stg4_s1[86 ]), .c(stg4_c1[86 ]), .co(stg4_co1[86 ]));
counter_5to3 u_a41_87 (.i0(stg3_s1_w[87 ]), .i1(stg3_c1_w[86 ]), .i2(stg3_s2_w[55 ]), .i3(stg3_c2_w[54 ]), .ci(stg4_co1[86 ]), .s(stg4_s1[87 ]), .c(stg4_c1[87 ]), .co(stg4_co1[87 ]));
counter_5to3 u_a41_88 (.i0(stg3_s1_w[88 ]), .i1(stg3_c1_w[87 ]), .i2(stg3_s2_w[56 ]), .i3(stg3_c2_w[55 ]), .ci(stg4_co1[87 ]), .s(stg4_s1[88 ]), .c(stg4_c1[88 ]), .co(stg4_co1[88 ]));
counter_5to3 u_a41_89 (.i0(stg3_s1_w[89 ]), .i1(stg3_c1_w[88 ]), .i2(stg3_s2_w[57 ]), .i3(stg3_c2_w[56 ]), .ci(stg4_co1[88 ]), .s(stg4_s1[89 ]), .c(stg4_c1[89 ]), .co(stg4_co1[89 ]));
counter_5to3 u_a41_90 (.i0(stg3_s1_w[90 ]), .i1(stg3_c1_w[89 ]), .i2(stg3_s2_w[58 ]), .i3(stg3_c2_w[57 ]), .ci(stg4_co1[89 ]), .s(stg4_s1[90 ]), .c(stg4_c1[90 ]), .co(stg4_co1[90 ]));
counter_5to3 u_a41_91 (.i0(stg3_s1_w[91 ]), .i1(stg3_c1_w[90 ]), .i2(stg3_s2_w[59 ]), .i3(stg3_c2_w[58 ]), .ci(stg4_co1[90 ]), .s(stg4_s1[91 ]), .c(stg4_c1[91 ]), .co(stg4_co1[91 ]));
counter_5to3 u_a41_92 (.i0(stg3_s1_w[92 ]), .i1(stg3_c1_w[91 ]), .i2(stg3_s2_w[60 ]), .i3(stg3_c2_w[59 ]), .ci(stg4_co1[91 ]), .s(stg4_s1[92 ]), .c(stg4_c1[92 ]), .co(stg4_co1[92 ]));
counter_5to3 u_a41_93 (.i0(stg3_s1_w[93 ]), .i1(stg3_c1_w[92 ]), .i2(stg3_s2_w[61 ]), .i3(stg3_c2_w[60 ]), .ci(stg4_co1[92 ]), .s(stg4_s1[93 ]), .c(stg4_c1[93 ]), .co(stg4_co1[93 ]));
counter_5to3 u_a41_94 (.i0(stg3_s1_w[94 ]), .i1(stg3_c1_w[93 ]), .i2(stg3_s2_w[62 ]), .i3(stg3_c2_w[61 ]), .ci(stg4_co1[93 ]), .s(stg4_s1[94 ]), .c(stg4_c1[94 ]), .co(stg4_co1[94 ]));
counter_5to3 u_a41_95 (.i0(stg3_s1_w[95 ]), .i1(stg3_c1_w[94 ]), .i2(stg3_s2_w[63 ]), .i3(stg3_c2_w[62 ]), .ci(stg4_co1[94 ]), .s(stg4_s1[95 ]), .c(stg4_c1[95 ]), .co(stg4_co1[95 ]));
counter_5to3 u_a41_96 (.i0(stg3_s1_w[96 ]), .i1(stg3_c1_w[95 ]), .i2(stg3_s2_w[64 ]), .i3(stg3_c2_w[63 ]), .ci(stg4_co1[95 ]), .s(stg4_s1[96 ]), .c(stg4_c1[96 ]), .co(stg4_co1[96 ]));
counter_5to3 u_a41_97 (.i0(stg3_s1_w[97 ]), .i1(stg3_c1_w[96 ]), .i2(stg3_s2_w[65 ]), .i3(stg3_c2_w[64 ]), .ci(stg4_co1[96 ]), .s(stg4_s1[97 ]), .c(stg4_c1[97 ]), .co(stg4_co1[97 ]));
counter_5to3 u_a41_98 (.i0(stg3_s1_w[98 ]), .i1(stg3_c1_w[97 ]), .i2(stg3_s2_w[66 ]), .i3(stg3_c2_w[65 ]), .ci(stg4_co1[97 ]), .s(stg4_s1[98 ]), .c(stg4_c1[98 ]), .co(stg4_co1[98 ]));
counter_5to3 u_a41_99 (.i0(stg3_s1_w[99 ]), .i1(stg3_c1_w[98 ]), .i2(stg3_s2_w[67 ]), .i3(stg3_c2_w[66 ]), .ci(stg4_co1[98 ]), .s(stg4_s1[99 ]), .c(stg4_c1[99 ]), .co(stg4_co1[99 ]));
counter_5to3 u_a41_100(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[99 ]), .i2(stg3_s2_w[68 ]), .i3(stg3_c2_w[67 ]), .ci(stg4_co1[99 ]), .s(stg4_s1[100]), .c(stg4_c1[100]), .co(stg4_co1[100]));
counter_5to3 u_a41_101(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[69 ]), .i3(stg3_c2_w[68 ]), .ci(stg4_co1[100]), .s(stg4_s1[101]), .c(stg4_c1[101]), .co(stg4_co1[101]));
counter_5to3 u_a41_102(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[70 ]), .i3(stg3_c2_w[69 ]), .ci(stg4_co1[101]), .s(stg4_s1[102]), .c(stg4_c1[102]), .co(stg4_co1[102]));
counter_5to3 u_a41_103(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[71 ]), .i3(stg3_c2_w[70 ]), .ci(stg4_co1[102]), .s(stg4_s1[103]), .c(stg4_c1[103]), .co(stg4_co1[103]));
counter_5to3 u_a41_104(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[72 ]), .i3(stg3_c2_w[71 ]), .ci(stg4_co1[103]), .s(stg4_s1[104]), .c(stg4_c1[104]), .co(stg4_co1[104]));
counter_5to3 u_a41_105(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[73 ]), .i3(stg3_c2_w[72 ]), .ci(stg4_co1[104]), .s(stg4_s1[105]), .c(stg4_c1[105]), .co(stg4_co1[105]));
counter_5to3 u_a41_106(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[74 ]), .i3(stg3_c2_w[73 ]), .ci(stg4_co1[105]), .s(stg4_s1[106]), .c(stg4_c1[106]), .co(stg4_co1[106]));
counter_5to3 u_a41_107(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[75 ]), .i3(stg3_c2_w[74 ]), .ci(stg4_co1[106]), .s(stg4_s1[107]), .c(stg4_c1[107]), .co(stg4_co1[107]));
counter_5to3 u_a41_108(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[76 ]), .i3(stg3_c2_w[75 ]), .ci(stg4_co1[107]), .s(stg4_s1[108]), .c(stg4_c1[108]), .co(stg4_co1[108]));
counter_5to3 u_a41_109(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[77 ]), .i3(stg3_c2_w[76 ]), .ci(stg4_co1[108]), .s(stg4_s1[109]), .c(stg4_c1[109]), .co(stg4_co1[109]));
counter_5to3 u_a41_110(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[78 ]), .i3(stg3_c2_w[77 ]), .ci(stg4_co1[109]), .s(stg4_s1[110]), .c(stg4_c1[110]), .co(stg4_co1[110]));
counter_5to3 u_a41_111(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[79 ]), .i3(stg3_c2_w[78 ]), .ci(stg4_co1[110]), .s(stg4_s1[111]), .c(stg4_c1[111]), .co(stg4_co1[111]));
counter_5to3 u_a41_112(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[80 ]), .i3(stg3_c2_w[79 ]), .ci(stg4_co1[111]), .s(stg4_s1[112]), .c(stg4_c1[112]), .co(stg4_co1[112]));
counter_5to3 u_a41_113(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[81 ]), .i3(stg3_c2_w[80 ]), .ci(stg4_co1[112]), .s(stg4_s1[113]), .c(stg4_c1[113]), .co(stg4_co1[113]));
counter_5to3 u_a41_114(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[82 ]), .i3(stg3_c2_w[81 ]), .ci(stg4_co1[113]), .s(stg4_s1[114]), .c(stg4_c1[114]), .co(stg4_co1[114]));
counter_5to3 u_a41_115(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[83 ]), .i3(stg3_c2_w[82 ]), .ci(stg4_co1[114]), .s(stg4_s1[115]), .c(stg4_c1[115]), .co(stg4_co1[115]));
counter_5to3 u_a41_116(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[84 ]), .i3(stg3_c2_w[83 ]), .ci(stg4_co1[115]), .s(stg4_s1[116]), .c(stg4_c1[116]), .co(stg4_co1[116]));
counter_5to3 u_a41_117(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[85 ]), .i3(stg3_c2_w[84 ]), .ci(stg4_co1[116]), .s(stg4_s1[117]), .c(stg4_c1[117]), .co(stg4_co1[117]));
counter_5to3 u_a41_118(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[86 ]), .i3(stg3_c2_w[85 ]), .ci(stg4_co1[117]), .s(stg4_s1[118]), .c(stg4_c1[118]), .co(stg4_co1[118]));
counter_5to3 u_a41_119(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[87 ]), .i3(stg3_c2_w[86 ]), .ci(stg4_co1[118]), .s(stg4_s1[119]), .c(stg4_c1[119]), .co(stg4_co1[119]));
counter_5to3 u_a41_120(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[88 ]), .i3(stg3_c2_w[87 ]), .ci(stg4_co1[119]), .s(stg4_s1[120]), .c(stg4_c1[120]), .co(stg4_co1[120]));
counter_5to3 u_a41_121(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[89 ]), .i3(stg3_c2_w[88 ]), .ci(stg4_co1[120]), .s(stg4_s1[121]), .c(stg4_c1[121]), .co(stg4_co1[121]));
counter_5to3 u_a41_122(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[90 ]), .i3(stg3_c2_w[89 ]), .ci(stg4_co1[121]), .s(stg4_s1[122]), .c(stg4_c1[122]), .co(stg4_co1[122]));
counter_5to3 u_a41_123(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[91 ]), .i3(stg3_c2_w[90 ]), .ci(stg4_co1[122]), .s(stg4_s1[123]), .c(stg4_c1[123]), .co(stg4_co1[123]));
counter_5to3 u_a41_124(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[92 ]), .i3(stg3_c2_w[91 ]), .ci(stg4_co1[123]), .s(stg4_s1[124]), .c(stg4_c1[124]), .co(stg4_co1[124]));
counter_5to3 u_a41_125(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[93 ]), .i3(stg3_c2_w[92 ]), .ci(stg4_co1[124]), .s(stg4_s1[125]), .c(stg4_c1[125]), .co(stg4_co1[125]));
counter_5to3 u_a41_126(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[94 ]), .i3(stg3_c2_w[93 ]), .ci(stg4_co1[125]), .s(stg4_s1[126]), .c(stg4_c1[126]), .co(stg4_co1[126]));
counter_5to3 u_a41_127(.i0(stg3_s1_w[100]), .i1(stg3_c1_w[100]), .i2(stg3_s2_w[95 ]), .i3(stg3_c2_w[94 ]), .ci(stg4_co1[126]), .s(stg4_s1[127]), .c(stg4_c1[127]), .co(stg4_co1[127]));

//================ fifth stage ================
wire [127:0] stg4_s1_w, stg4_c1_w;
wire [65:0]  pp33_w4;

// ========= pipeline ==============
reg [127:0] stg4_s1_ff, stg4_c1_ff;
reg [65:0]  pp33_f4;

always @(posedge clk or negedge rstn)begin
    if(!rstn)begin
        stg4_s1_ff <= 128'b0;
        stg4_c1_ff <= 128'b0;
        pp33_f4    <= 66'b0;
    end
    else begin
        stg4_s1_ff <= stg4_s1;
        stg4_c1_ff <= stg4_c1;
        pp33_f4    <= pp33_w3;
    end
end

assign stg4_s1_w   = stg4_s1_ff;
assign stg4_c1_w   = stg4_c1_ff;
assign pp33_w4     = pp33_f4   ;

wire [127:0] stg5_s1, stg5_c1, stg5_co1;

// =========================== fifth stage 1st group ============================================================================================================
assign stg5_s1[0]  = stg4_s1_w[0];
assign stg5_co1[0] = 1'b0;
half_adder u_a51_0  (.a(stg4_s1_w[1  ]), .b(stg4_c1_w[0  ]), .s(stg5_s1[1  ]), .co(stg5_co1[1 ]));
half_adder u_a51_1  (.a(stg4_s1_w[2  ]), .b(stg4_c1_w[1  ]), .s(stg5_s1[2  ]), .co(stg5_co1[2 ]));
half_adder u_a51_2  (.a(stg4_s1_w[3  ]), .b(stg4_c1_w[2  ]), .s(stg5_s1[3  ]), .co(stg5_co1[3 ]));
half_adder u_a51_3  (.a(stg4_s1_w[4  ]), .b(stg4_c1_w[3  ]), .s(stg5_s1[4  ]), .co(stg5_co1[4 ]));
half_adder u_a51_4  (.a(stg4_s1_w[5  ]), .b(stg4_c1_w[4  ]), .s(stg5_s1[5  ]), .co(stg5_co1[5 ]));
half_adder u_a51_5  (.a(stg4_s1_w[6  ]), .b(stg4_c1_w[5  ]), .s(stg5_s1[6  ]), .co(stg5_co1[6 ]));
half_adder u_a51_6  (.a(stg4_s1_w[7  ]), .b(stg4_c1_w[6  ]), .s(stg5_s1[7  ]), .co(stg5_co1[7 ]));
half_adder u_a51_7  (.a(stg4_s1_w[8  ]), .b(stg4_c1_w[7  ]), .s(stg5_s1[8  ]), .co(stg5_co1[8 ]));
half_adder u_a51_8  (.a(stg4_s1_w[9  ]), .b(stg4_c1_w[8  ]), .s(stg5_s1[9  ]), .co(stg5_co1[9 ]));
half_adder u_a51_9  (.a(stg4_s1_w[10 ]), .b(stg4_c1_w[9  ]), .s(stg5_s1[10 ]), .co(stg5_co1[10]));
half_adder u_a51_10 (.a(stg4_s1_w[11 ]), .b(stg4_c1_w[10 ]), .s(stg5_s1[11 ]), .co(stg5_co1[11]));
half_adder u_a51_11 (.a(stg4_s1_w[12 ]), .b(stg4_c1_w[11 ]), .s(stg5_s1[12 ]), .co(stg5_co1[12]));
half_adder u_a51_12 (.a(stg4_s1_w[13 ]), .b(stg4_c1_w[12 ]), .s(stg5_s1[13 ]), .co(stg5_co1[13]));
half_adder u_a51_13 (.a(stg4_s1_w[14 ]), .b(stg4_c1_w[13 ]), .s(stg5_s1[14 ]), .co(stg5_co1[14]));
half_adder u_a51_14 (.a(stg4_s1_w[15 ]), .b(stg4_c1_w[14 ]), .s(stg5_s1[15 ]), .co(stg5_co1[15]));
half_adder u_a51_15 (.a(stg4_s1_w[16 ]), .b(stg4_c1_w[15 ]), .s(stg5_s1[16 ]), .co(stg5_co1[16]));
half_adder u_a51_16 (.a(stg4_s1_w[17 ]), .b(stg4_c1_w[16 ]), .s(stg5_s1[17 ]), .co(stg5_co1[17]));
half_adder u_a51_17 (.a(stg4_s1_w[18 ]), .b(stg4_c1_w[17 ]), .s(stg5_s1[18 ]), .co(stg5_co1[18]));
half_adder u_a51_18 (.a(stg4_s1_w[19 ]), .b(stg4_c1_w[18 ]), .s(stg5_s1[19 ]), .co(stg5_co1[19]));
half_adder u_a51_19 (.a(stg4_s1_w[20 ]), .b(stg4_c1_w[19 ]), .s(stg5_s1[20 ]), .co(stg5_co1[20]));
half_adder u_a51_20 (.a(stg4_s1_w[21 ]), .b(stg4_c1_w[20 ]), .s(stg5_s1[21 ]), .co(stg5_co1[21]));
half_adder u_a51_21 (.a(stg4_s1_w[22 ]), .b(stg4_c1_w[21 ]), .s(stg5_s1[22 ]), .co(stg5_co1[22]));
half_adder u_a51_22 (.a(stg4_s1_w[23 ]), .b(stg4_c1_w[22 ]), .s(stg5_s1[23 ]), .co(stg5_co1[23]));
half_adder u_a51_23 (.a(stg4_s1_w[24 ]), .b(stg4_c1_w[23 ]), .s(stg5_s1[24 ]), .co(stg5_co1[24]));
half_adder u_a51_24 (.a(stg4_s1_w[25 ]), .b(stg4_c1_w[24 ]), .s(stg5_s1[25 ]), .co(stg5_co1[25]));
half_adder u_a51_25 (.a(stg4_s1_w[26 ]), .b(stg4_c1_w[25 ]), .s(stg5_s1[26 ]), .co(stg5_co1[26]));
half_adder u_a51_26 (.a(stg4_s1_w[27 ]), .b(stg4_c1_w[26 ]), .s(stg5_s1[27 ]), .co(stg5_co1[27]));
half_adder u_a51_27 (.a(stg4_s1_w[28 ]), .b(stg4_c1_w[27 ]), .s(stg5_s1[28 ]), .co(stg5_co1[28]));
half_adder u_a51_28 (.a(stg4_s1_w[29 ]), .b(stg4_c1_w[28 ]), .s(stg5_s1[29 ]), .co(stg5_co1[29]));
half_adder u_a51_29 (.a(stg4_s1_w[30 ]), .b(stg4_c1_w[29 ]), .s(stg5_s1[30 ]), .co(stg5_co1[30]));
half_adder u_a51_30 (.a(stg4_s1_w[31 ]), .b(stg4_c1_w[30 ]), .s(stg5_s1[31 ]), .co(stg5_co1[31]));
half_adder u_a51_31 (.a(stg4_s1_w[32 ]), .b(stg4_c1_w[31 ]), .s(stg5_s1[32 ]), .co(stg5_co1[32]));
half_adder u_a51_32 (.a(stg4_s1_w[33 ]), .b(stg4_c1_w[32 ]), .s(stg5_s1[33 ]), .co(stg5_co1[33]));
half_adder u_a51_33 (.a(stg4_s1_w[34 ]), .b(stg4_c1_w[33 ]), .s(stg5_s1[34 ]), .co(stg5_co1[34]));
half_adder u_a51_34 (.a(stg4_s1_w[35 ]), .b(stg4_c1_w[34 ]), .s(stg5_s1[35 ]), .co(stg5_co1[35]));
half_adder u_a51_35 (.a(stg4_s1_w[36 ]), .b(stg4_c1_w[35 ]), .s(stg5_s1[36 ]), .co(stg5_co1[36]));
half_adder u_a51_36 (.a(stg4_s1_w[37 ]), .b(stg4_c1_w[36 ]), .s(stg5_s1[37 ]), .co(stg5_co1[37]));
half_adder u_a51_37 (.a(stg4_s1_w[38 ]), .b(stg4_c1_w[37 ]), .s(stg5_s1[38 ]), .co(stg5_co1[38]));
half_adder u_a51_38 (.a(stg4_s1_w[39 ]), .b(stg4_c1_w[38 ]), .s(stg5_s1[39 ]), .co(stg5_co1[39]));
half_adder u_a51_39 (.a(stg4_s1_w[40 ]), .b(stg4_c1_w[39 ]), .s(stg5_s1[40 ]), .co(stg5_co1[40]));
half_adder u_a51_40 (.a(stg4_s1_w[41 ]), .b(stg4_c1_w[40 ]), .s(stg5_s1[41 ]), .co(stg5_co1[41]));
half_adder u_a51_41 (.a(stg4_s1_w[42 ]), .b(stg4_c1_w[41 ]), .s(stg5_s1[42 ]), .co(stg5_co1[42]));
half_adder u_a51_42 (.a(stg4_s1_w[43 ]), .b(stg4_c1_w[42 ]), .s(stg5_s1[43 ]), .co(stg5_co1[43]));
half_adder u_a51_43 (.a(stg4_s1_w[44 ]), .b(stg4_c1_w[43 ]), .s(stg5_s1[44 ]), .co(stg5_co1[44]));
half_adder u_a51_44 (.a(stg4_s1_w[45 ]), .b(stg4_c1_w[44 ]), .s(stg5_s1[45 ]), .co(stg5_co1[45]));
half_adder u_a51_45 (.a(stg4_s1_w[46 ]), .b(stg4_c1_w[45 ]), .s(stg5_s1[46 ]), .co(stg5_co1[46]));
half_adder u_a51_46 (.a(stg4_s1_w[47 ]), .b(stg4_c1_w[46 ]), .s(stg5_s1[47 ]), .co(stg5_co1[47]));
half_adder u_a51_47 (.a(stg4_s1_w[48 ]), .b(stg4_c1_w[47 ]), .s(stg5_s1[48 ]), .co(stg5_co1[48]));
half_adder u_a51_48 (.a(stg4_s1_w[49 ]), .b(stg4_c1_w[48 ]), .s(stg5_s1[49 ]), .co(stg5_co1[49]));
half_adder u_a51_49 (.a(stg4_s1_w[50 ]), .b(stg4_c1_w[49 ]), .s(stg5_s1[50 ]), .co(stg5_co1[50]));
half_adder u_a51_50 (.a(stg4_s1_w[51 ]), .b(stg4_c1_w[50 ]), .s(stg5_s1[51 ]), .co(stg5_co1[51]));
half_adder u_a51_51 (.a(stg4_s1_w[52 ]), .b(stg4_c1_w[51 ]), .s(stg5_s1[52 ]), .co(stg5_co1[52]));
half_adder u_a51_52 (.a(stg4_s1_w[53 ]), .b(stg4_c1_w[52 ]), .s(stg5_s1[53 ]), .co(stg5_co1[53]));
half_adder u_a51_53 (.a(stg4_s1_w[54 ]), .b(stg4_c1_w[53 ]), .s(stg5_s1[54 ]), .co(stg5_co1[54]));
half_adder u_a51_54 (.a(stg4_s1_w[55 ]), .b(stg4_c1_w[54 ]), .s(stg5_s1[55 ]), .co(stg5_co1[55]));
half_adder u_a51_55 (.a(stg4_s1_w[56 ]), .b(stg4_c1_w[55 ]), .s(stg5_s1[56 ]), .co(stg5_co1[56]));
half_adder u_a51_56 (.a(stg4_s1_w[57 ]), .b(stg4_c1_w[56 ]), .s(stg5_s1[57 ]), .co(stg5_co1[57]));
half_adder u_a51_57 (.a(stg4_s1_w[58 ]), .b(stg4_c1_w[57 ]), .s(stg5_s1[58 ]), .co(stg5_co1[58]));
half_adder u_a51_58 (.a(stg4_s1_w[59 ]), .b(stg4_c1_w[58 ]), .s(stg5_s1[59 ]), .co(stg5_co1[59]));
half_adder u_a51_59 (.a(stg4_s1_w[60 ]), .b(stg4_c1_w[59 ]), .s(stg5_s1[60 ]), .co(stg5_co1[60]));
half_adder u_a51_60 (.a(stg4_s1_w[61 ]), .b(stg4_c1_w[60 ]), .s(stg5_s1[61 ]), .co(stg5_co1[61]));
half_adder u_a51_61 (.a(stg4_s1_w[62 ]), .b(stg4_c1_w[61 ]), .s(stg5_s1[62 ]), .co(stg5_co1[62]));
half_adder u_a51_62 (.a(stg4_s1_w[63 ]), .b(stg4_c1_w[62 ]), .s(stg5_s1[63 ]), .co(stg5_co1[63]));

full_adder u_a51_63 (.a(stg4_s1_w[64 ]), .b(stg4_c1_w[63 ]), .ci(pp33_w4[0 ]  ), .s(stg5_s1[64 ]), .co(stg5_co1[64 ]));
full_adder u_a51_64 (.a(stg4_s1_w[65 ]), .b(stg4_c1_w[64 ]), .ci(pp33_w4[1 ]  ), .s(stg5_s1[65 ]), .co(stg5_co1[65 ]));
full_adder u_a51_65 (.a(stg4_s1_w[66 ]), .b(stg4_c1_w[65 ]), .ci(pp33_w4[2 ]  ), .s(stg5_s1[66 ]), .co(stg5_co1[66 ]));
full_adder u_a51_66 (.a(stg4_s1_w[67 ]), .b(stg4_c1_w[66 ]), .ci(pp33_w4[3 ]  ), .s(stg5_s1[67 ]), .co(stg5_co1[67 ]));
full_adder u_a51_67 (.a(stg4_s1_w[68 ]), .b(stg4_c1_w[67 ]), .ci(pp33_w4[4 ]  ), .s(stg5_s1[68 ]), .co(stg5_co1[68 ]));
full_adder u_a51_68 (.a(stg4_s1_w[69 ]), .b(stg4_c1_w[68 ]), .ci(pp33_w4[5 ]  ), .s(stg5_s1[69 ]), .co(stg5_co1[69 ]));
full_adder u_a51_69 (.a(stg4_s1_w[70 ]), .b(stg4_c1_w[69 ]), .ci(pp33_w4[6 ]  ), .s(stg5_s1[70 ]), .co(stg5_co1[70 ]));
full_adder u_a51_70 (.a(stg4_s1_w[71 ]), .b(stg4_c1_w[70 ]), .ci(pp33_w4[7 ]  ), .s(stg5_s1[71 ]), .co(stg5_co1[71 ]));
full_adder u_a51_71 (.a(stg4_s1_w[72 ]), .b(stg4_c1_w[71 ]), .ci(pp33_w4[8 ]  ), .s(stg5_s1[72 ]), .co(stg5_co1[72 ]));
full_adder u_a51_72 (.a(stg4_s1_w[73 ]), .b(stg4_c1_w[72 ]), .ci(pp33_w4[9 ]  ), .s(stg5_s1[73 ]), .co(stg5_co1[73 ]));
full_adder u_a51_73 (.a(stg4_s1_w[74 ]), .b(stg4_c1_w[73 ]), .ci(pp33_w4[10]  ), .s(stg5_s1[74 ]), .co(stg5_co1[74 ]));
full_adder u_a51_74 (.a(stg4_s1_w[75 ]), .b(stg4_c1_w[74 ]), .ci(pp33_w4[11]  ), .s(stg5_s1[75 ]), .co(stg5_co1[75 ]));
full_adder u_a51_75 (.a(stg4_s1_w[76 ]), .b(stg4_c1_w[75 ]), .ci(pp33_w4[12]  ), .s(stg5_s1[76 ]), .co(stg5_co1[76 ]));
full_adder u_a51_76 (.a(stg4_s1_w[77 ]), .b(stg4_c1_w[76 ]), .ci(pp33_w4[13]  ), .s(stg5_s1[77 ]), .co(stg5_co1[77 ]));
full_adder u_a51_77 (.a(stg4_s1_w[78 ]), .b(stg4_c1_w[77 ]), .ci(pp33_w4[14]  ), .s(stg5_s1[78 ]), .co(stg5_co1[78 ]));
full_adder u_a51_78 (.a(stg4_s1_w[79 ]), .b(stg4_c1_w[78 ]), .ci(pp33_w4[15]  ), .s(stg5_s1[79 ]), .co(stg5_co1[79 ]));
full_adder u_a51_79 (.a(stg4_s1_w[80 ]), .b(stg4_c1_w[79 ]), .ci(pp33_w4[16]  ), .s(stg5_s1[80 ]), .co(stg5_co1[80 ]));
full_adder u_a51_80 (.a(stg4_s1_w[81 ]), .b(stg4_c1_w[80 ]), .ci(pp33_w4[17]  ), .s(stg5_s1[81 ]), .co(stg5_co1[81 ]));
full_adder u_a51_81 (.a(stg4_s1_w[82 ]), .b(stg4_c1_w[81 ]), .ci(pp33_w4[18]  ), .s(stg5_s1[82 ]), .co(stg5_co1[82 ]));
full_adder u_a51_82 (.a(stg4_s1_w[83 ]), .b(stg4_c1_w[82 ]), .ci(pp33_w4[19]  ), .s(stg5_s1[83 ]), .co(stg5_co1[83 ]));
full_adder u_a51_83 (.a(stg4_s1_w[84 ]), .b(stg4_c1_w[83 ]), .ci(pp33_w4[20]  ), .s(stg5_s1[84 ]), .co(stg5_co1[84 ]));
full_adder u_a51_84 (.a(stg4_s1_w[85 ]), .b(stg4_c1_w[84 ]), .ci(pp33_w4[21]  ), .s(stg5_s1[85 ]), .co(stg5_co1[85 ]));
full_adder u_a51_85 (.a(stg4_s1_w[86 ]), .b(stg4_c1_w[85 ]), .ci(pp33_w4[22]  ), .s(stg5_s1[86 ]), .co(stg5_co1[86 ]));
full_adder u_a51_86 (.a(stg4_s1_w[87 ]), .b(stg4_c1_w[86 ]), .ci(pp33_w4[23]  ), .s(stg5_s1[87 ]), .co(stg5_co1[87 ]));
full_adder u_a51_87 (.a(stg4_s1_w[88 ]), .b(stg4_c1_w[87 ]), .ci(pp33_w4[24]  ), .s(stg5_s1[88 ]), .co(stg5_co1[88 ]));
full_adder u_a51_88 (.a(stg4_s1_w[89 ]), .b(stg4_c1_w[88 ]), .ci(pp33_w4[25]  ), .s(stg5_s1[89 ]), .co(stg5_co1[89 ]));
full_adder u_a51_89 (.a(stg4_s1_w[90 ]), .b(stg4_c1_w[89 ]), .ci(pp33_w4[26]  ), .s(stg5_s1[90 ]), .co(stg5_co1[90 ]));
full_adder u_a51_90 (.a(stg4_s1_w[91 ]), .b(stg4_c1_w[90 ]), .ci(pp33_w4[27]  ), .s(stg5_s1[91 ]), .co(stg5_co1[91 ]));
full_adder u_a51_91 (.a(stg4_s1_w[92 ]), .b(stg4_c1_w[91 ]), .ci(pp33_w4[28]  ), .s(stg5_s1[92 ]), .co(stg5_co1[92 ]));
full_adder u_a51_92 (.a(stg4_s1_w[93 ]), .b(stg4_c1_w[92 ]), .ci(pp33_w4[29]  ), .s(stg5_s1[93 ]), .co(stg5_co1[93 ]));
full_adder u_a51_93 (.a(stg4_s1_w[94 ]), .b(stg4_c1_w[93 ]), .ci(pp33_w4[30]  ), .s(stg5_s1[94 ]), .co(stg5_co1[94 ]));
full_adder u_a51_94 (.a(stg4_s1_w[95 ]), .b(stg4_c1_w[94 ]), .ci(pp33_w4[31]  ), .s(stg5_s1[95 ]), .co(stg5_co1[95 ]));
full_adder u_a51_95 (.a(stg4_s1_w[96 ]), .b(stg4_c1_w[95 ]), .ci(pp33_w4[32]  ), .s(stg5_s1[96 ]), .co(stg5_co1[96 ]));
full_adder u_a51_96 (.a(stg4_s1_w[97 ]), .b(stg4_c1_w[96 ]), .ci(pp33_w4[33]  ), .s(stg5_s1[97 ]), .co(stg5_co1[97 ]));
full_adder u_a51_97 (.a(stg4_s1_w[98 ]), .b(stg4_c1_w[97 ]), .ci(pp33_w4[34]  ), .s(stg5_s1[98 ]), .co(stg5_co1[98 ]));
full_adder u_a51_98 (.a(stg4_s1_w[99 ]), .b(stg4_c1_w[98 ]), .ci(pp33_w4[35]  ), .s(stg5_s1[99 ]), .co(stg5_co1[99 ]));
full_adder u_a51_99 (.a(stg4_s1_w[100]), .b(stg4_c1_w[99 ]), .ci(pp33_w4[36]  ), .s(stg5_s1[100]), .co(stg5_co1[100]));
full_adder u_a51_100(.a(stg4_s1_w[101]), .b(stg4_c1_w[100]), .ci(pp33_w4[37]  ), .s(stg5_s1[101]), .co(stg5_co1[101]));
full_adder u_a51_101(.a(stg4_s1_w[102]), .b(stg4_c1_w[101]), .ci(pp33_w4[38]  ), .s(stg5_s1[102]), .co(stg5_co1[102]));
full_adder u_a51_102(.a(stg4_s1_w[103]), .b(stg4_c1_w[102]), .ci(pp33_w4[39]  ), .s(stg5_s1[103]), .co(stg5_co1[103]));
full_adder u_a51_103(.a(stg4_s1_w[104]), .b(stg4_c1_w[103]), .ci(pp33_w4[40]  ), .s(stg5_s1[104]), .co(stg5_co1[104]));
full_adder u_a51_104(.a(stg4_s1_w[105]), .b(stg4_c1_w[104]), .ci(pp33_w4[41]  ), .s(stg5_s1[105]), .co(stg5_co1[105]));
full_adder u_a51_105(.a(stg4_s1_w[106]), .b(stg4_c1_w[105]), .ci(pp33_w4[42]  ), .s(stg5_s1[106]), .co(stg5_co1[106]));
full_adder u_a51_106(.a(stg4_s1_w[107]), .b(stg4_c1_w[106]), .ci(pp33_w4[43]  ), .s(stg5_s1[107]), .co(stg5_co1[107]));
full_adder u_a51_107(.a(stg4_s1_w[108]), .b(stg4_c1_w[107]), .ci(pp33_w4[44]  ), .s(stg5_s1[108]), .co(stg5_co1[108]));
full_adder u_a51_108(.a(stg4_s1_w[109]), .b(stg4_c1_w[108]), .ci(pp33_w4[45]  ), .s(stg5_s1[109]), .co(stg5_co1[109]));
full_adder u_a51_109(.a(stg4_s1_w[110]), .b(stg4_c1_w[109]), .ci(pp33_w4[46]  ), .s(stg5_s1[110]), .co(stg5_co1[110]));
full_adder u_a51_110(.a(stg4_s1_w[111]), .b(stg4_c1_w[110]), .ci(pp33_w4[47]  ), .s(stg5_s1[111]), .co(stg5_co1[111]));
full_adder u_a51_111(.a(stg4_s1_w[112]), .b(stg4_c1_w[111]), .ci(pp33_w4[48]  ), .s(stg5_s1[112]), .co(stg5_co1[112]));
full_adder u_a51_112(.a(stg4_s1_w[113]), .b(stg4_c1_w[112]), .ci(pp33_w4[49]  ), .s(stg5_s1[113]), .co(stg5_co1[113]));
full_adder u_a51_113(.a(stg4_s1_w[114]), .b(stg4_c1_w[113]), .ci(pp33_w4[50]  ), .s(stg5_s1[114]), .co(stg5_co1[114]));
full_adder u_a51_114(.a(stg4_s1_w[115]), .b(stg4_c1_w[114]), .ci(pp33_w4[51]  ), .s(stg5_s1[115]), .co(stg5_co1[115]));
full_adder u_a51_115(.a(stg4_s1_w[116]), .b(stg4_c1_w[115]), .ci(pp33_w4[52]  ), .s(stg5_s1[116]), .co(stg5_co1[116]));
full_adder u_a51_116(.a(stg4_s1_w[117]), .b(stg4_c1_w[116]), .ci(pp33_w4[53]  ), .s(stg5_s1[117]), .co(stg5_co1[117]));
full_adder u_a51_117(.a(stg4_s1_w[118]), .b(stg4_c1_w[117]), .ci(pp33_w4[54]  ), .s(stg5_s1[118]), .co(stg5_co1[118]));
full_adder u_a51_118(.a(stg4_s1_w[119]), .b(stg4_c1_w[118]), .ci(pp33_w4[55]  ), .s(stg5_s1[119]), .co(stg5_co1[119]));
full_adder u_a51_119(.a(stg4_s1_w[120]), .b(stg4_c1_w[119]), .ci(pp33_w4[56]  ), .s(stg5_s1[120]), .co(stg5_co1[120]));
full_adder u_a51_120(.a(stg4_s1_w[121]), .b(stg4_c1_w[120]), .ci(pp33_w4[57]  ), .s(stg5_s1[121]), .co(stg5_co1[121]));
full_adder u_a51_121(.a(stg4_s1_w[122]), .b(stg4_c1_w[121]), .ci(pp33_w4[58]  ), .s(stg5_s1[122]), .co(stg5_co1[122]));
full_adder u_a51_122(.a(stg4_s1_w[123]), .b(stg4_c1_w[122]), .ci(pp33_w4[59]  ), .s(stg5_s1[123]), .co(stg5_co1[123]));
full_adder u_a51_123(.a(stg4_s1_w[124]), .b(stg4_c1_w[123]), .ci(pp33_w4[60]  ), .s(stg5_s1[124]), .co(stg5_co1[124]));
full_adder u_a51_124(.a(stg4_s1_w[125]), .b(stg4_c1_w[124]), .ci(pp33_w4[61]  ), .s(stg5_s1[125]), .co(stg5_co1[125]));
full_adder u_a51_125(.a(stg4_s1_w[126]), .b(stg4_c1_w[125]), .ci(pp33_w4[62]  ), .s(stg5_s1[126]), .co(stg5_co1[126]));
full_adder u_a51_126(.a(stg4_s1_w[127]), .b(stg4_c1_w[126]), .ci(pp33_w4[63]  ), .s(stg5_s1[127]), .co(stg5_co1[127]));

// ================== final result ===================

wire [127:0] stg5_s1_w, stg5_co1_w;

// ============== pipeline ================
reg [127:0] stg5_s1_ff, stg5_co1_ff;

always @(posedge clk or negedge rstn)begin
    if (!rstn)begin
        stg5_s1_ff  <= 0;
        stg5_co1_ff <= 0;
    end
    else begin
        stg5_s1_ff  <= stg5_s1;
        stg5_co1_ff <= stg5_co1;
    end
end

assign stg5_s1_w = stg5_s1_ff;
assign stg5_co1_w = stg5_co1_ff;

assign final_p = stg5_s1_w + {stg5_co1_w[126:0], 1'b0};

endmodule
